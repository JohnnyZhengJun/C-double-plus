VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO A2O1A1I_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN A2O1A1I_xp33_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.144 0.728 0.288 0.8 ;
        RECT 0.216 0.28 0.288 0.8 ;
        RECT 0.14 0.28 0.288 0.352 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.728 0.576 0.8 ;
        RECT 0.504 0.28 0.576 0.8 ;
        RECT 0.428 0.28 0.576 0.352 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.868 0.352 ;
        RECT 0.72 0.688 0.864 0.76 ;
        RECT 0.72 0.28 0.792 0.76 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.08 0.688 1.224 0.76 ;
        RECT 1.152 0.3 1.224 0.76 ;
        RECT 1.048 0.3 1.224 0.372 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.856 0.86 1.44 0.932 ;
        RECT 1.368 0.148 1.44 0.932 ;
        RECT 1.24 0.148 1.44 0.22 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.116 0.18 ;
      RECT 0.16 0.9 0.704 0.972 ;
  END
END A2O1A1I_xp33_75t

MACRO A2O1A1O1I_xp25_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN A2O1A1O1I_xp25_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.504 0.576 0.576 ;
        RECT 0.36 0.756 0.508 0.828 ;
        RECT 0.36 0.252 0.508 0.324 ;
        RECT 0.36 0.252 0.432 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.14 0.756 0.288 0.828 ;
        RECT 0.216 0.252 0.288 0.828 ;
        RECT 0.14 0.252 0.288 0.324 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.756 0.792 0.828 ;
        RECT 0.72 0.252 0.792 0.828 ;
        RECT 0.644 0.252 0.792 0.324 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.756 1.084 0.828 ;
        RECT 0.936 0.252 1.084 0.324 ;
        RECT 0.936 0.252 1.008 0.828 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.508 1.676 0.58 ;
        RECT 1.368 0.756 1.516 0.828 ;
        RECT 1.368 0.252 1.516 0.324 ;
        RECT 1.368 0.252 1.44 0.828 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.692 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.044 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.828 0.9 1.548 0.972 ;
      RECT 0.16 0.108 0.9 0.18 ;
      RECT 0.16 0.9 0.684 0.972 ;
  END
END A2O1A1O1I_xp25_75t

MACRO AND2_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_x1_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.312 0.504 0.8 ;
        RECT 0.356 0.312 0.504 0.384 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.668 0.308 0.74 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.312 0.22 0.384 ;
        RECT 0.072 0.312 0.144 0.972 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.808 0.108 1.008 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.684 0.972 ;
      RECT 0.612 0.648 0.684 0.972 ;
      RECT 0.612 0.648 0.792 0.72 ;
      RECT 0.72 0.396 0.792 0.72 ;
      RECT 0.612 0.396 0.792 0.468 ;
      RECT 0.612 0.16 0.684 0.468 ;
      RECT 0.26 0.16 0.684 0.232 ;
  END
END AND2_x1_75t

MACRO AND2_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_x2_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.356 0.728 0.576 0.8 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.136 0.144 0.972 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.828 0.108 1.224 0.18 ;
        RECT 0.828 0.736 0.9 0.972 ;
        RECT 0.828 0.108 0.9 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.72 0.972 ;
      RECT 0.648 0.108 0.72 0.972 ;
      RECT 0.648 0.504 0.812 0.576 ;
      RECT 0.28 0.108 0.352 0.344 ;
      RECT 0.28 0.108 0.72 0.18 ;
  END
END AND2_x2_75t

MACRO AND2_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_x4_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.112 1.008 0.6 ;
        RECT 0.072 0.112 1.008 0.184 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.112 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.9 0.576 0.972 ;
        RECT 0.504 0.428 0.576 0.972 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.24 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.72 0.9 0.924 0.972 ;
      RECT 0.72 0.256 0.792 0.972 ;
      RECT 0.72 0.728 1.224 0.8 ;
      RECT 1.152 0.484 1.224 0.8 ;
      RECT 0.46 0.256 0.792 0.328 ;
  END
END AND2_x4_75t

MACRO AND2_x6_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_x6_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.112 1.008 0.6 ;
        RECT 0.072 0.112 1.008 0.184 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.112 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.728 0.576 0.8 ;
        RECT 0.504 0.428 0.576 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 2.216 0.972 ;
        RECT 1.24 0.108 2.216 0.18 ;
        RECT 1.8 0.108 1.872 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.924 0.972 ;
      RECT 0.72 0.256 0.792 0.972 ;
      RECT 0.72 0.728 1.224 0.8 ;
      RECT 1.152 0.484 1.224 0.8 ;
      RECT 0.46 0.256 0.792 0.328 ;
  END
END AND2_x6_75t

MACRO AND3_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_x1_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.14 0.756 0.288 0.828 ;
        RECT 0.216 0.252 0.288 0.828 ;
        RECT 0.14 0.252 0.288 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.504 0.576 0.576 ;
        RECT 0.36 0.728 0.504 0.8 ;
        RECT 0.36 0.28 0.504 0.352 ;
        RECT 0.36 0.28 0.432 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.756 0.792 0.828 ;
        RECT 0.72 0.28 0.792 0.828 ;
        RECT 0.648 0.28 0.792 0.352 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.732 1.224 0.804 ;
        RECT 1.152 0.304 1.224 0.804 ;
        RECT 1.044 0.304 1.224 0.376 ;
        RECT 1.044 0.732 1.116 0.94 ;
        RECT 1.044 0.136 1.116 0.376 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.936 0.972 ;
      RECT 0.864 0.108 0.936 0.972 ;
      RECT 0.864 0.504 1.052 0.576 ;
      RECT 0.16 0.108 0.936 0.18 ;
  END
END AND3_x1_75t

MACRO AND3_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_x2_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.14 0.756 0.288 0.828 ;
        RECT 0.216 0.252 0.288 0.828 ;
        RECT 0.14 0.252 0.288 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.504 0.576 0.576 ;
        RECT 0.36 0.756 0.508 0.828 ;
        RECT 0.36 0.252 0.508 0.324 ;
        RECT 0.36 0.252 0.432 0.828 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.756 0.792 0.828 ;
        RECT 0.72 0.252 0.792 0.828 ;
        RECT 0.644 0.252 0.792 0.324 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.044 0.108 1.44 0.18 ;
        RECT 1.044 0.736 1.116 0.972 ;
        RECT 1.044 0.108 1.116 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.936 0.972 ;
      RECT 0.864 0.108 0.936 0.972 ;
      RECT 0.864 0.504 1.136 0.576 ;
      RECT 0.16 0.108 0.936 0.18 ;
  END
END AND3_x2_75t

MACRO AND3_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_x4_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.756 2.812 0.828 ;
        RECT 2.448 0.396 2.812 0.468 ;
        RECT 2.448 0.396 2.52 0.828 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.756 2.348 0.828 ;
        RECT 2.016 0.396 2.348 0.468 ;
        RECT 2.016 0.396 2.088 0.828 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.728 1.516 0.8 ;
        RECT 1.368 0.28 1.516 0.352 ;
        RECT 1.368 0.28 1.44 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.92 0.972 ;
        RECT 0.072 0.108 0.92 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.04 0.9 2.984 0.972 ;
      RECT 2.912 0.108 2.984 0.972 ;
      RECT 1.04 0.168 1.112 0.972 ;
      RECT 0.872 0.504 1.112 0.576 ;
      RECT 2.536 0.108 2.984 0.18 ;
      RECT 1.888 0.252 2.804 0.324 ;
      RECT 1.24 0.108 2.216 0.18 ;
  END
END AND3_x4_75t

MACRO AND3_x6_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_x6_75t 0 0 ;
  SIZE 3.456 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.808 0.504 3.104 0.576 ;
        RECT 2.808 0.748 2.956 0.82 ;
        RECT 2.808 0.432 2.88 0.82 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.504 2.54 0.576 ;
        RECT 2.232 0.748 2.38 0.82 ;
        RECT 2.232 0.448 2.304 0.82 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.724 0.748 1.872 0.82 ;
        RECT 1.8 0.26 1.872 0.82 ;
        RECT 1.672 0.504 1.872 0.576 ;
        RECT 1.724 0.26 1.872 0.332 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.456 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.9 1.352 0.972 ;
        RECT 0.18 0.108 1.352 0.18 ;
        RECT 0.18 0.108 0.252 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.476 0.9 3.384 0.972 ;
      RECT 3.312 0.28 3.384 0.972 ;
      RECT 1.476 0.504 1.548 0.972 ;
      RECT 1.348 0.504 1.548 0.576 ;
      RECT 2.968 0.28 3.384 0.352 ;
      RECT 2.016 0.252 2.648 0.324 ;
      RECT 2.016 0.108 2.088 0.324 ;
      RECT 1.672 0.108 2.088 0.18 ;
      RECT 2.32 0.108 3.296 0.18 ;
  END
END AND3_x6_75t

MACRO AND4_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4_x1_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.28 0.364 0.352 ;
        RECT 0.216 0.28 0.288 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.728 0.576 0.8 ;
        RECT 0.504 0.256 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.108 0.792 0.8 ;
        RECT 0.644 0.108 0.792 0.18 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.136 1.008 0.656 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.196 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.24 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 1.008 0.972 ;
      RECT 0.936 0.756 1.008 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.936 0.756 1.224 0.828 ;
      RECT 1.152 0.48 1.224 0.828 ;
      RECT 0.072 0.108 0.34 0.18 ;
  END
END AND4_x1_75t

MACRO AND4_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4_x2_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.252 0.364 0.324 ;
        RECT 0.216 0.252 0.288 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.388 0.756 0.576 0.828 ;
        RECT 0.504 0.256 0.576 0.828 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.108 0.792 0.8 ;
        RECT 0.644 0.108 0.792 0.18 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.656 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.196 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.24 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 1.008 0.972 ;
      RECT 0.936 0.756 1.008 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.936 0.756 1.224 0.828 ;
      RECT 1.152 0.464 1.224 0.828 ;
      RECT 0.072 0.108 0.292 0.18 ;
  END
END AND4_x2_75t

MACRO AND4_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4_x4_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.26 0.364 0.332 ;
        RECT 0.216 0.26 0.288 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.388 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.108 0.792 0.8 ;
        RECT 0.644 0.108 0.792 0.18 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.656 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.196 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.24 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 1.008 0.972 ;
      RECT 0.936 0.756 1.008 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.936 0.756 1.224 0.828 ;
      RECT 1.152 0.464 1.224 0.828 ;
      RECT 0.072 0.108 0.292 0.18 ;
  END
END AND4_x4_75t

MACRO AND4_x6_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4_x6_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.26 0.364 0.332 ;
        RECT 0.216 0.26 0.288 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.388 0.756 0.576 0.828 ;
        RECT 0.504 0.26 0.576 0.828 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.108 0.792 0.8 ;
        RECT 0.644 0.108 0.792 0.18 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.136 1.008 0.656 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.196 0.9 2.304 0.972 ;
        RECT 2.232 0.108 2.304 0.972 ;
        RECT 1.24 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 1.008 0.972 ;
      RECT 0.936 0.756 1.008 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.936 0.756 1.224 0.828 ;
      RECT 1.152 0.464 1.224 0.828 ;
      RECT 0.072 0.108 0.292 0.18 ;
  END
END AND4_x6_75t

MACRO AND5_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND5_x1_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.756 0.364 0.828 ;
        RECT 0.216 0.252 0.364 0.324 ;
        RECT 0.216 0.252 0.288 0.828 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.256 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.108 0.792 0.8 ;
        RECT 0.644 0.108 0.792 0.18 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.256 1.008 0.8 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.108 1.224 0.656 ;
        RECT 1.076 0.108 1.224 0.18 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.396 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 1.4 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 1.224 0.972 ;
      RECT 1.152 0.756 1.224 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 1.152 0.756 1.44 0.828 ;
      RECT 1.368 0.464 1.44 0.828 ;
      RECT 0.072 0.108 0.292 0.18 ;
  END
END AND5_x1_75t

MACRO AND5_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND5_x2_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.956 0.552 2.028 0.8 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.684 1.008 0.756 ;
        RECT 0.936 0.252 1.008 0.756 ;
        RECT 0.808 0.252 1.008 0.324 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.708 0.576 2.54 0.648 ;
      LAYER M1 ;
        RECT 2.448 0.484 2.52 0.668 ;
        RECT 1.728 0.556 1.8 0.74 ;
      LAYER V1 ;
        RECT 1.728 0.576 1.8 0.648 ;
        RECT 2.448 0.576 2.52 0.648 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.564 0.432 2.756 0.504 ;
      LAYER M1 ;
        RECT 2.664 0.412 2.736 0.592 ;
        RECT 1.584 0.412 1.656 0.592 ;
      LAYER V1 ;
        RECT 1.584 0.432 1.656 0.504 ;
        RECT 2.664 0.432 2.736 0.504 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.268 0.576 1.46 0.648 ;
      LAYER M1 ;
        RECT 1.368 0.452 1.44 0.668 ;
        RECT 0.288 0.552 0.36 0.812 ;
      LAYER V1 ;
        RECT 0.288 0.576 0.36 0.648 ;
        RECT 1.368 0.576 1.44 0.648 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.42 0.432 1.244 0.504 ;
      LAYER M1 ;
        RECT 1.152 0.412 1.224 0.592 ;
        RECT 0.44 0.412 0.512 0.592 ;
      LAYER V1 ;
        RECT 0.44 0.432 0.512 0.504 ;
        RECT 1.152 0.432 1.224 0.504 ;
    END
  END E
  OBS
    LAYER M1 ;
      RECT 2.772 0.144 2.844 0.308 ;
      RECT 2.752 0.144 2.9 0.216 ;
      RECT 0.612 0.9 2.864 0.972 ;
      RECT 2.124 0.34 2.196 0.972 ;
      RECT 0.612 0.504 0.684 0.972 ;
      RECT 0.612 0.504 0.812 0.576 ;
      RECT 2.556 0.108 2.628 0.308 ;
      RECT 1.692 0.108 1.764 0.308 ;
      RECT 1.692 0.108 2.628 0.18 ;
      RECT 1.476 0.144 1.548 0.308 ;
      RECT 1.436 0.144 1.584 0.216 ;
      RECT 1.26 0.108 1.332 0.308 ;
      RECT 0.396 0.108 0.468 0.272 ;
      RECT 0.396 0.108 1.332 0.18 ;
      RECT 0.18 0.144 0.252 0.376 ;
      RECT 0.124 0.144 0.272 0.216 ;
      RECT 2.32 0.288 2.432 0.36 ;
      RECT 1.888 0.288 2 0.36 ;
    LAYER M2 ;
      RECT 0.16 0.144 2.864 0.216 ;
      RECT 1.852 0.288 2.432 0.36 ;
    LAYER V1 ;
      RECT 2.772 0.144 2.844 0.216 ;
      RECT 2.34 0.288 2.412 0.36 ;
      RECT 1.908 0.288 1.98 0.36 ;
      RECT 1.476 0.144 1.548 0.216 ;
      RECT 0.18 0.144 0.252 0.216 ;
  END
END AND5_x2_75t

MACRO AO211_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO211_x2_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.588 0.728 2.736 0.8 ;
        RECT 2.664 0.28 2.736 0.8 ;
        RECT 2.588 0.28 2.736 0.352 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.576 0.576 0.648 ;
        RECT 0.504 0.256 0.576 0.648 ;
        RECT 0.072 0.576 0.144 0.776 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.888 0.728 2.088 0.8 ;
        RECT 2.016 0.28 2.088 0.8 ;
        RECT 1.888 0.28 2.088 0.352 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.492 0.432 2.324 0.504 ;
      LAYER M1 ;
        RECT 2.232 0.412 2.304 0.596 ;
        RECT 1.512 0.412 1.584 0.596 ;
      LAYER V1 ;
        RECT 1.512 0.432 1.584 0.504 ;
        RECT 2.232 0.432 2.304 0.504 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.052 0.288 1.028 0.36 ;
      LAYER M1 ;
        RECT 0.916 0.288 1.028 0.36 ;
        RECT 0.936 0.288 1.008 0.488 ;
        RECT 0.072 0.2 0.316 0.272 ;
        RECT 0.072 0.2 0.144 0.38 ;
      LAYER V1 ;
        RECT 0.072 0.288 0.144 0.36 ;
        RECT 0.936 0.288 1.008 0.36 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.648 0.108 0.72 0.756 ;
      RECT 1.692 0.504 1.892 0.576 ;
      RECT 1.692 0.108 1.764 0.576 ;
      RECT 0.648 0.108 2.648 0.18 ;
      RECT 0.828 0.72 1.028 0.792 ;
      RECT 0.828 0.628 0.9 0.792 ;
      RECT 0.16 0.9 2.864 0.972 ;
      RECT 0.268 0.72 0.488 0.792 ;
    LAYER M2 ;
      RECT 0.268 0.72 1.028 0.792 ;
    LAYER V1 ;
      RECT 0.92 0.72 0.992 0.792 ;
      RECT 0.288 0.72 0.36 0.792 ;
  END
END AO211_x2_75t

MACRO AO21_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21_x1_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.076 0.756 1.224 0.828 ;
        RECT 1.152 0.136 1.224 0.828 ;
        RECT 0.916 0.504 1.224 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.26 0.868 0.332 ;
        RECT 0.72 0.26 0.792 0.656 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.332 0.972 ;
        RECT 0.072 0.152 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.216 0.756 0.92 0.828 ;
      RECT 0.216 0.108 0.288 0.828 ;
      RECT 0.216 0.108 0.704 0.18 ;
      RECT 0.592 0.9 1.136 0.972 ;
  END
END AO21_x1_75t

MACRO AO21_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21_x2_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.136 0.144 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.792 0.28 0.864 0.656 ;
        RECT 0.7 0.504 0.864 0.576 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.92 0.9 1.44 0.972 ;
        RECT 1.368 0.276 1.44 0.972 ;
        RECT 1.08 0.276 1.44 0.348 ;
        RECT 1.08 0.152 1.152 0.348 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.756 1.008 0.828 ;
      RECT 0.936 0.108 1.008 0.828 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.16 0.9 0.704 0.972 ;
  END
END AO21_x2_75t

MACRO AO221_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221_x1_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.084 0.352 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.252 1.44 0.632 ;
        RECT 1.204 0.504 1.44 0.576 ;
        RECT 1.292 0.252 1.44 0.324 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.28 0.364 0.352 ;
        RECT 0.216 0.28 0.288 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.584 0.576 0.656 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.888 0.9 2.088 0.972 ;
        RECT 2.016 0.108 2.088 0.972 ;
        RECT 1.836 0.108 2.088 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.756 0.504 0.828 ;
      RECT 0.072 0.108 0.144 0.828 ;
      RECT 1.584 0.504 1.896 0.576 ;
      RECT 1.584 0.108 1.656 0.576 ;
      RECT 0.072 0.108 1.656 0.18 ;
      RECT 0.8 0.756 1.356 0.828 ;
      RECT 0.156 0.9 0.704 0.972 ;
  END
END AO221_x1_75t

MACRO AO221_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO221_x2_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.26 1.084 0.332 ;
        RECT 0.936 0.26 1.008 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.26 1.44 0.676 ;
        RECT 1.204 0.504 1.44 0.576 ;
        RECT 1.292 0.26 1.44 0.332 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.26 0.364 0.332 ;
        RECT 0.216 0.26 0.288 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.604 0.576 0.676 ;
        RECT 0.504 0.392 0.576 0.676 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.26 0.792 0.656 ;
        RECT 0.644 0.26 0.792 0.332 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.888 0.9 2.196 0.972 ;
        RECT 2.124 0.108 2.196 0.972 ;
        RECT 1.836 0.108 2.196 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.756 0.504 0.828 ;
      RECT 0.072 0.108 0.144 0.828 ;
      RECT 1.584 0.504 1.896 0.576 ;
      RECT 1.584 0.108 1.656 0.576 ;
      RECT 0.072 0.108 1.656 0.18 ;
      RECT 0.8 0.756 1.356 0.828 ;
      RECT 0.156 0.9 0.704 0.972 ;
  END
END AO221_x2_75t

MACRO AO222_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222_x1_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.316 0.792 0.596 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.316 0.576 0.596 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.316 2.088 0.62 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.316 1.872 0.62 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.304 0.316 1.376 0.62 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.316 1.656 0.64 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.72 0.272 0.792 ;
        RECT 0.144 0.224 0.216 0.432 ;
        RECT 0.072 0.36 0.144 0.792 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.72 1.568 0.792 ;
      RECT 1.044 0.144 1.116 0.792 ;
      RECT 0.268 0.504 0.432 0.576 ;
      RECT 0.36 0.144 0.432 0.576 ;
      RECT 0.36 0.144 2.216 0.216 ;
      RECT 2.104 0.864 2.252 0.936 ;
      RECT 1.908 0.7 1.98 0.848 ;
      RECT 1.636 0.864 1.784 0.936 ;
      RECT 1.204 0.864 1.352 0.936 ;
      RECT 0.592 0.72 0.704 0.792 ;
    LAYER M2 ;
      RECT 1.24 0.864 2.216 0.936 ;
      RECT 0.592 0.72 2 0.792 ;
    LAYER V1 ;
      RECT 2.124 0.864 2.196 0.936 ;
      RECT 1.908 0.72 1.98 0.792 ;
      RECT 1.692 0.864 1.764 0.936 ;
      RECT 1.26 0.864 1.332 0.936 ;
      RECT 0.612 0.72 0.684 0.792 ;
  END
END AO222_x1_75t

MACRO AO222_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO222_x2_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.512 0.28 1.584 0.688 ;
        RECT 1.436 0.28 1.584 0.352 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.728 1.948 0.8 ;
        RECT 1.8 0.28 1.872 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.612 1.084 0.684 ;
        RECT 0.936 0.26 1.084 0.332 ;
        RECT 0.936 0.26 1.008 0.684 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.504 0.812 0.576 ;
        RECT 0.648 0.28 0.72 0.648 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.612 0.364 0.684 ;
        RECT 0.216 0.252 0.364 0.324 ;
        RECT 0.216 0.252 0.288 0.684 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.648 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.104 0.9 2.52 0.972 ;
        RECT 2.448 0.108 2.52 0.972 ;
        RECT 2.124 0.108 2.52 0.18 ;
        RECT 2.124 0.108 2.196 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.756 0.488 0.828 ;
      RECT 0.072 0.108 0.144 0.828 ;
      RECT 1.944 0.504 2.216 0.576 ;
      RECT 1.944 0.108 2.016 0.576 ;
      RECT 0.072 0.108 2.016 0.18 ;
      RECT 1.368 0.9 1.872 0.972 ;
      RECT 1.368 0.756 1.44 0.972 ;
      RECT 0.808 0.756 1.44 0.828 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END AO222_x2_75t

MACRO AO22_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22_x1_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.392 0.576 0.828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.26 1.084 0.332 ;
        RECT 0.936 0.26 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.26 0.792 0.656 ;
        RECT 0.644 0.26 0.792 0.332 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.672 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.756 1.44 0.828 ;
      RECT 1.368 0.108 1.44 0.828 ;
      RECT 1.368 0.504 1.676 0.576 ;
      RECT 0.592 0.108 1.44 0.18 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END AO22_x1_75t

MACRO AO22_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22_x2_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.424 0.728 0.576 0.8 ;
        RECT 0.504 0.392 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.084 0.324 ;
        RECT 0.936 0.252 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.26 0.792 0.656 ;
        RECT 0.644 0.26 0.792 0.332 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.9 2.088 0.972 ;
        RECT 2.016 0.108 2.088 0.972 ;
        RECT 1.672 0.108 2.088 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.756 1.44 0.828 ;
      RECT 1.368 0.108 1.44 0.828 ;
      RECT 1.368 0.504 1.676 0.576 ;
      RECT 0.428 0.108 1.44 0.18 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END AO22_x2_75t

MACRO AO31_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31_x1_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.284 0.576 0.688 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.108 0.792 0.8 ;
        RECT 0.644 0.108 0.792 0.18 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.8 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.748 0.436 0.82 ;
        RECT 0.288 0.28 0.36 0.82 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.24 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.144 0.668 0.216 0.876 ;
      RECT 0.072 0.108 0.144 0.74 ;
      RECT 0.072 0.108 0.488 0.18 ;
      RECT 1.152 0.28 1.224 0.716 ;
      RECT 0.376 0.9 0.92 0.972 ;
    LAYER M2 ;
      RECT 0.052 0.576 1.244 0.648 ;
    LAYER V1 ;
      RECT 1.152 0.576 1.224 0.648 ;
      RECT 0.072 0.576 0.144 0.648 ;
  END
END AO31_x1_75t

MACRO AO31_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO31_x2_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.584 0.828 ;
        RECT 0.512 0.304 0.584 0.828 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.728 0.728 2.876 0.8 ;
        RECT 2.728 0.108 2.876 0.18 ;
        RECT 2.728 0.108 2.8 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.512 0.304 1.584 0.776 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.836 0.72 2.144 0.792 ;
        RECT 0.204 0.432 2.108 0.504 ;
      LAYER M1 ;
        RECT 1.996 0.72 2.144 0.792 ;
        RECT 2.016 0.412 2.088 0.792 ;
        RECT 0.836 0.508 1.044 0.58 ;
        RECT 0.836 0.72 0.984 0.792 ;
        RECT 0.836 0.508 0.908 0.792 ;
        RECT 0.224 0.304 0.296 0.6 ;
      LAYER V1 ;
        RECT 0.224 0.432 0.296 0.504 ;
        RECT 0.892 0.72 0.964 0.792 ;
        RECT 2.016 0.72 2.088 0.792 ;
        RECT 2.016 0.432 2.088 0.504 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.132 0.288 1.892 0.36 ;
      LAYER M1 ;
        RECT 1.78 0.288 1.892 0.36 ;
        RECT 1.8 0.288 1.872 0.6 ;
        RECT 1.152 0.28 1.224 0.6 ;
      LAYER V1 ;
        RECT 1.152 0.288 1.224 0.36 ;
        RECT 1.8 0.288 1.872 0.36 ;
    END
  END A3
  OBS
    LAYER M1 ;
      RECT 2.34 0.276 2.412 0.668 ;
      RECT 2.34 0.276 2.628 0.348 ;
      RECT 2.556 0.16 2.628 0.348 ;
      RECT 0.16 0.9 2.864 0.972 ;
      RECT 2.556 0.556 2.628 0.74 ;
      RECT 0.16 0.108 2 0.18 ;
      RECT 1.368 0.476 1.44 0.668 ;
      RECT 0.856 0.288 0.968 0.36 ;
      RECT 0.656 0.304 0.728 0.668 ;
      RECT 0.368 0.28 0.44 0.468 ;
    LAYER M2 ;
      RECT 0.636 0.576 2.648 0.648 ;
      RECT 0.348 0.288 0.968 0.36 ;
    LAYER V1 ;
      RECT 2.556 0.576 2.628 0.648 ;
      RECT 2.34 0.576 2.412 0.648 ;
      RECT 1.368 0.576 1.44 0.648 ;
      RECT 0.876 0.288 0.948 0.36 ;
      RECT 0.656 0.576 0.728 0.648 ;
      RECT 0.368 0.288 0.44 0.36 ;
  END
END AO31_x2_75t

MACRO AO322_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO322_x2_75t 0 0 ;
  SIZE 3.24 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.612 1.3 0.684 ;
        RECT 1.152 0.252 1.3 0.324 ;
        RECT 1.152 0.252 1.224 0.684 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.252 2.164 0.324 ;
        RECT 2.016 0.252 2.088 0.656 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.24 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.536 0.9 3.168 0.972 ;
        RECT 3.096 0.108 3.168 0.972 ;
        RECT 2.536 0.108 3.168 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.584 0.756 2.304 0.828 ;
      RECT 2.232 0.504 2.304 0.828 ;
      RECT 1.584 0.108 1.656 0.828 ;
      RECT 2.232 0.504 2.972 0.576 ;
      RECT 0.16 0.108 1.784 0.18 ;
      RECT 0.376 0.9 0.792 0.972 ;
      RECT 0.72 0.756 0.792 0.972 ;
      RECT 0.72 0.756 1.352 0.828 ;
      RECT 1.024 0.9 2 0.972 ;
  END
END AO322_x2_75t

MACRO AO32_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32_x1_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.392 1.008 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.756 0.792 0.828 ;
        RECT 0.72 0.28 0.792 0.828 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.688 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.252 1.224 0.656 ;
        RECT 1.076 0.252 1.224 0.324 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.252 0.252 0.324 ;
        RECT 0.18 0.136 0.252 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.24 0.756 1.656 0.828 ;
      RECT 1.584 0.108 1.656 0.828 ;
      RECT 0.26 0.504 0.432 0.576 ;
      RECT 0.36 0.108 0.432 0.576 ;
      RECT 0.36 0.108 1.656 0.18 ;
      RECT 0.592 0.9 1.568 0.972 ;
  END
END AO32_x1_75t

MACRO AO32_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO32_x2_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.756 1.32 0.828 ;
        RECT 1.152 0.28 1.224 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.728 0.792 0.8 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.656 0.28 1.728 0.656 ;
        RECT 1.58 0.28 1.728 0.352 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.488 0.972 ;
        RECT 0.072 0.272 0.468 0.344 ;
        RECT 0.396 0.148 0.468 0.344 ;
        RECT 0.072 0.272 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.456 0.756 1.872 0.828 ;
      RECT 1.8 0.108 1.872 0.828 ;
      RECT 0.372 0.504 0.648 0.576 ;
      RECT 0.576 0.108 0.648 0.576 ;
      RECT 0.576 0.108 1.872 0.18 ;
      RECT 0.808 0.9 1.784 0.972 ;
  END
END AO32_x2_75t

MACRO AO331_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO331_x1_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.324 0.18 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.884 0.9 2.088 0.972 ;
      RECT 2.016 0.108 2.088 0.972 ;
      RECT 0.288 0.252 0.36 0.608 ;
      RECT 0.288 0.252 0.576 0.324 ;
      RECT 0.504 0.108 0.576 0.324 ;
      RECT 0.504 0.108 2.088 0.18 ;
      RECT 1.232 0.756 1.788 0.828 ;
      RECT 0.584 0.9 1.572 0.972 ;
  END
END AO331_x1_75t

MACRO AO331_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO331_x2_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END B3
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.28 2.088 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.108 0.54 0.18 ;
        RECT 0.288 0.9 0.488 0.972 ;
        RECT 0.288 0.108 0.36 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.1 0.9 2.304 0.972 ;
      RECT 2.232 0.108 2.304 0.972 ;
      RECT 0.504 0.252 0.576 0.608 ;
      RECT 0.504 0.252 0.792 0.324 ;
      RECT 0.72 0.108 0.792 0.324 ;
      RECT 0.72 0.108 2.304 0.18 ;
      RECT 1.448 0.756 2.004 0.828 ;
      RECT 0.8 0.9 1.788 0.972 ;
  END
END AO331_x2_75t

MACRO AO332_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO332_x1_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.28 2.088 0.656 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.376 0.18 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.884 0.756 2.304 0.828 ;
      RECT 2.232 0.108 2.304 0.828 ;
      RECT 0.288 0.252 0.36 0.604 ;
      RECT 0.288 0.252 0.576 0.324 ;
      RECT 0.504 0.108 0.576 0.324 ;
      RECT 0.504 0.108 2.304 0.18 ;
      RECT 0.584 0.9 1.008 0.972 ;
      RECT 0.936 0.756 1.008 0.972 ;
      RECT 0.936 0.756 1.572 0.828 ;
      RECT 1.232 0.9 2.224 0.972 ;
  END
END AO332_x1_75t

MACRO AO332_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO332_x2_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.28 2.304 0.656 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.28 2.088 0.656 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.592 0.18 ;
        RECT 0.072 0.9 0.488 0.972 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.1 0.756 2.52 0.828 ;
      RECT 2.448 0.108 2.52 0.828 ;
      RECT 0.504 0.252 0.576 0.604 ;
      RECT 0.504 0.252 0.792 0.324 ;
      RECT 0.72 0.108 0.792 0.324 ;
      RECT 0.72 0.108 2.52 0.18 ;
      RECT 0.8 0.9 1.224 0.972 ;
      RECT 1.152 0.756 1.224 0.972 ;
      RECT 1.152 0.756 1.788 0.828 ;
      RECT 1.448 0.9 2.44 0.972 ;
  END
END AO332_x2_75t

MACRO AO333_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO333_x1_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.656 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.28 2.304 0.656 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.28 2.088 0.656 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.324 0.18 ;
        RECT 0.072 0.9 0.276 0.972 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.884 0.9 2.52 0.972 ;
      RECT 2.448 0.108 2.52 0.972 ;
      RECT 0.288 0.252 0.36 0.608 ;
      RECT 0.288 0.252 0.576 0.324 ;
      RECT 0.504 0.108 0.576 0.324 ;
      RECT 0.504 0.108 2.52 0.18 ;
      RECT 1.24 0.756 2.304 0.828 ;
      RECT 0.592 0.9 1.58 0.972 ;
  END
END AO333_x1_75t

MACRO AO333_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO333_x2_75t 0 0 ;
  SIZE 2.808 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.28 2.52 0.656 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.28 2.304 0.656 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.28 2.088 0.656 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.808 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.488 0.972 ;
        RECT 0.072 0.324 0.468 0.396 ;
        RECT 0.396 0.18 0.468 0.396 ;
        RECT 0.072 0.324 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.1 0.9 2.736 0.972 ;
      RECT 2.664 0.108 2.736 0.972 ;
      RECT 0.268 0.504 0.648 0.576 ;
      RECT 0.576 0.108 0.648 0.576 ;
      RECT 0.576 0.108 2.736 0.18 ;
      RECT 1.456 0.756 2.52 0.828 ;
      RECT 0.808 0.9 1.796 0.972 ;
  END
END AO333_x2_75t

MACRO AO33_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO33_x1_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.392 1.008 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.26 0.792 0.8 ;
        RECT 0.644 0.26 0.792 0.332 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.728 0.576 0.8 ;
        RECT 0.504 0.392 0.576 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.26 1.224 0.632 ;
        RECT 1.076 0.26 1.224 0.332 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.304 1.44 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.656 0.28 1.728 0.656 ;
        RECT 1.58 0.28 1.728 0.352 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.144 0.34 0.216 0.72 ;
        RECT 0.072 0.648 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.24 0.756 1.872 0.828 ;
      RECT 1.8 0.108 1.872 0.828 ;
      RECT 0.288 0.108 0.36 0.596 ;
      RECT 0.288 0.108 1.872 0.18 ;
      RECT 0.592 0.9 1.568 0.972 ;
  END
END AO33_x1_75t

MACRO AO33_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO33_x2_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.748 1.3 0.82 ;
        RECT 1.152 0.28 1.224 0.82 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.728 0.792 0.8 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.488 0.972 ;
        RECT 0.072 0.272 0.468 0.344 ;
        RECT 0.396 0.148 0.468 0.344 ;
        RECT 0.072 0.272 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.456 0.756 2.088 0.828 ;
      RECT 2.016 0.108 2.088 0.828 ;
      RECT 0.268 0.504 0.648 0.576 ;
      RECT 0.576 0.108 0.648 0.576 ;
      RECT 0.576 0.108 2.088 0.18 ;
      RECT 0.796 0.9 1.796 0.972 ;
  END
END AO33_x2_75t

MACRO AOI211_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211_x1_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.72 0.748 1.872 0.82 ;
        RECT 1.8 0.108 1.872 0.82 ;
        RECT 1.72 0.108 1.872 0.18 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.748 1.52 0.82 ;
        RECT 1.368 0.304 1.52 0.376 ;
        RECT 1.368 0.304 1.44 0.82 ;
    END
  END A2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.304 0.684 0.608 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.204 0.288 1.028 0.36 ;
      LAYER M1 ;
        RECT 0.88 0.288 1.028 0.36 ;
        RECT 0.224 0.268 0.296 0.596 ;
      LAYER V1 ;
        RECT 0.224 0.288 0.296 0.36 ;
        RECT 0.936 0.288 1.008 0.36 ;
    END
  END B
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.584 0.72 1.148 0.792 ;
      LAYER M1 ;
        RECT 0.376 0.108 1.352 0.18 ;
        RECT 1.036 0.72 1.224 0.792 ;
        RECT 1.152 0.108 1.224 0.792 ;
        RECT 0.584 0.72 0.732 0.792 ;
      LAYER V1 ;
        RECT 0.612 0.72 0.684 0.792 ;
        RECT 1.056 0.72 1.128 0.792 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 2 0.972 ;
      RECT 0.84 0.556 0.912 0.74 ;
      RECT 0.396 0.556 0.468 0.74 ;
    LAYER M2 ;
      RECT 0.376 0.576 0.932 0.648 ;
    LAYER V1 ;
      RECT 0.84 0.576 0.912 0.648 ;
      RECT 0.396 0.576 0.468 0.648 ;
  END
END AOI211_x1_75t

MACRO AOI211_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211_xp5_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.612 0.576 0.684 ;
        RECT 0.504 0.392 0.576 0.684 ;
        RECT 0.428 0.392 0.576 0.464 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.26 0.792 0.656 ;
        RECT 0.644 0.26 0.792 0.332 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.16 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.704 0.972 ;
  END
END AOI211_xp5_75t

MACRO AOI21_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_x1_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 0.612 1.008 0.684 ;
        RECT 0.936 0.252 1.008 0.684 ;
        RECT 0.86 0.252 1.008 0.324 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.756 1.44 0.828 ;
        RECT 1.368 0.484 1.44 0.828 ;
        RECT 0.288 0.484 0.36 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.476 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.072 0.108 1.656 0.18 ;
        RECT 0.072 0.9 0.252 0.972 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.484 0.432 1.244 0.504 ;
      LAYER M1 ;
        RECT 1.152 0.412 1.224 0.596 ;
        RECT 0.504 0.412 0.576 0.596 ;
      LAYER V1 ;
        RECT 0.504 0.432 0.576 0.504 ;
        RECT 1.152 0.432 1.224 0.504 ;
    END
  END A1
  OBS
    LAYER M1 ;
      RECT 0.396 0.9 1.332 0.972 ;
  END
END AOI21_x1_75t

MACRO AOI21_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_xp33_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.5 0.38 0.572 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.716 0.728 0.864 0.8 ;
        RECT 0.792 0.26 0.864 0.8 ;
        RECT 0.716 0.26 0.864 0.332 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.428 0.108 1.008 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.684 0.972 ;
  END
END AOI21_xp33_75t

MACRO AOI21_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_xp5_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.728 0.576 0.8 ;
        RECT 0.504 0.28 0.576 0.8 ;
        RECT 0.428 0.28 0.576 0.352 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.5 0.38 0.572 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.716 0.728 0.864 0.8 ;
        RECT 0.792 0.28 0.864 0.8 ;
        RECT 0.716 0.28 0.864 0.352 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.568 0.108 1.008 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.684 0.972 ;
  END
END AOI21_xp5_75t

MACRO AOI221_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221_x1_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.612 0.868 0.684 ;
        RECT 0.72 0.108 0.792 0.684 ;
        RECT 0.644 0.108 0.792 0.18 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.324 1.3 0.396 ;
        RECT 1.076 0.612 1.224 0.684 ;
        RECT 1.152 0.324 1.224 0.684 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.612 1.948 0.684 ;
        RECT 1.8 0.324 1.872 0.684 ;
        RECT 1.564 0.504 1.872 0.576 ;
        RECT 1.724 0.324 1.872 0.396 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.504 2.544 0.576 ;
        RECT 2.156 0.756 2.304 0.828 ;
        RECT 2.232 0.324 2.304 0.828 ;
        RECT 2.156 0.324 2.304 0.396 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.536 0.756 2.952 0.828 ;
        RECT 2.88 0.18 2.952 0.828 ;
        RECT 1.024 0.18 2.952 0.252 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.008 0.972 ;
      RECT 0.936 0.756 1.008 0.972 ;
      RECT 0.936 0.756 2 0.828 ;
      RECT 1.24 0.9 2.864 0.972 ;
  END
END AOI221_x1_75t

MACRO AOI221_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221_xp5_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.136 1.224 0.656 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.92 0.18 ;
        RECT 0.072 0.756 0.492 0.828 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.804 0.756 1.356 0.828 ;
      RECT 0.16 0.9 0.704 0.972 ;
  END
END AOI221_xp5_75t

MACRO AOI222_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222_xp33_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.136 1.872 0.8 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 1.596 0.18 ;
        RECT 0.072 0.756 0.488 0.828 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.368 0.9 1.872 0.972 ;
      RECT 1.368 0.756 1.44 0.972 ;
      RECT 0.808 0.756 1.44 0.828 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END AOI222_xp33_75t

MACRO AOI22_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_x1_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.612 1.516 0.684 ;
        RECT 1.368 0.396 1.516 0.468 ;
        RECT 1.368 0.396 1.44 0.684 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.252 1.872 0.596 ;
        RECT 1.152 0.252 1.872 0.324 ;
        RECT 1.152 0.252 1.224 0.608 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.644 0.756 0.792 0.828 ;
        RECT 0.72 0.396 0.792 0.828 ;
        RECT 0.644 0.396 0.792 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.616 ;
        RECT 0.288 0.252 1.008 0.324 ;
        RECT 0.288 0.756 0.436 0.828 ;
        RECT 0.288 0.252 0.36 0.828 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.236 0.756 2.088 0.828 ;
        RECT 2.016 0.108 2.088 0.828 ;
        RECT 0.152 0.108 2.088 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 2 0.972 ;
  END
END AOI22_x1_75t

MACRO AOI22_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_xp33_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.504 0.596 0.576 ;
        RECT 0.432 0.756 0.58 0.828 ;
        RECT 0.432 0.256 0.504 0.828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.26 0.792 0.656 ;
        RECT 0.644 0.26 0.792 0.332 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.592 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END AOI22_xp33_75t

MACRO AOI22_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_xp5_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.26 0.576 0.828 ;
        RECT 0.428 0.26 0.576 0.332 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.592 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END AOI22_xp5_75t

MACRO AOI311_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI311_xp33_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.108 0.576 0.828 ;
        RECT 0.428 0.108 0.576 0.18 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 0.792 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.936 0.972 ;
  END
END AOI311_xp33_75t

MACRO AOI31_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31_xp33_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.26 0.792 0.8 ;
        RECT 0.644 0.26 0.792 0.34 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.432 0.5 0.596 0.572 ;
        RECT 0.432 0.748 0.58 0.82 ;
        RECT 0.432 0.108 0.58 0.18 ;
        RECT 0.432 0.108 0.504 0.82 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.804 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.372 0.9 0.92 0.972 ;
  END
END AOI31_xp33_75t

MACRO AOI31_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31_xp67_75t 0 0 ;
  SIZE 2.808 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.664 0.28 2.736 0.8 ;
        RECT 2.212 0.504 2.736 0.576 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.504 1.676 0.576 ;
        RECT 1.152 0.252 1.3 0.324 ;
        RECT 1.152 0.252 1.224 0.656 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.236 0.828 ;
        RECT 0.072 0.108 0.236 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 0.812 0.576 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.808 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.34 0.9 2.652 0.972 ;
        RECT 2.34 0.756 2.412 0.972 ;
        RECT 0.808 0.756 2.412 0.828 ;
        RECT 0.936 0.252 1.008 0.828 ;
        RECT 0.808 0.252 1.008 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 2.104 0.108 2.652 0.18 ;
      RECT 1.456 0.324 2.432 0.396 ;
      RECT 0.16 0.9 2.216 0.972 ;
      RECT 0.376 0.108 1.788 0.18 ;
  END
END AOI31_xp67_75t

MACRO AOI321_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI321_xp33_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.108 0.576 0.656 ;
        RECT 0.428 0.108 0.576 0.18 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.756 1.656 0.828 ;
        RECT 1.584 0.108 1.656 0.828 ;
        RECT 0.792 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.024 0.9 1.584 0.972 ;
      RECT 0.376 0.756 0.92 0.828 ;
  END
END AOI321_xp33_75t

MACRO AOI322_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI322_xp5_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.66 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.136 0.36 0.656 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.66 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.756 1.872 0.828 ;
        RECT 1.8 0.108 1.872 0.828 ;
        RECT 0.588 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.9 1.8 0.972 ;
      RECT 0.156 0.756 1.136 0.828 ;
  END
END AOI322_xp5_75t

MACRO AOI32_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32_x1_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.076 0.756 1.224 0.828 ;
        RECT 1.152 0.34 1.224 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.108 1.44 0.8 ;
        RECT 1.292 0.108 1.44 0.18 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.728 1.732 0.8 ;
        RECT 1.584 0.108 1.732 0.18 ;
        RECT 1.584 0.108 1.656 0.8 ;
    END
  END A3
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.612 0.668 0.684 ;
        RECT 0.504 0.252 0.652 0.324 ;
        RECT 0.504 0.252 0.576 0.684 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.052 0.144 1.156 0.216 ;
      LAYER M1 ;
        RECT 1.044 0.144 1.156 0.216 ;
        RECT 0.072 0.756 0.92 0.828 ;
        RECT 0.052 0.144 0.252 0.216 ;
        RECT 0.072 0.144 0.144 0.828 ;
      LAYER V1 ;
        RECT 0.072 0.144 0.144 0.216 ;
        RECT 1.064 0.144 1.136 0.216 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.268 0.432 1.028 0.504 ;
      LAYER M1 ;
        RECT 0.936 0.412 1.008 0.596 ;
        RECT 0.288 0.412 0.36 0.596 ;
      LAYER V1 ;
        RECT 0.288 0.432 0.36 0.504 ;
        RECT 0.936 0.432 1.008 0.504 ;
    END
  END B1
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.568 0.972 ;
      RECT 0.376 0.108 0.92 0.18 ;
  END
END AOI32_x1_75t

MACRO AOI32_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32_xp33_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.232 0.972 ;
        RECT 0.072 0.252 0.232 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.416 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.416 0.252 0.576 0.324 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.756 0.888 0.828 ;
        RECT 0.72 0.28 0.792 0.828 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.148 0.612 1.296 0.684 ;
        RECT 1.224 0.252 1.296 0.684 ;
        RECT 1.148 0.252 1.296 0.324 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.756 1.44 0.828 ;
        RECT 1.368 0.108 1.44 0.828 ;
        RECT 0.16 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 1.352 0.972 ;
  END
END AOI32_xp33_75t

MACRO AOI32_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32_xp67_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.076 0.756 1.224 0.828 ;
        RECT 1.152 0.34 1.224 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.108 1.44 0.8 ;
        RECT 1.292 0.108 1.44 0.18 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.728 1.732 0.8 ;
        RECT 1.584 0.108 1.732 0.18 ;
        RECT 1.584 0.108 1.656 0.8 ;
    END
  END A3
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.612 0.668 0.684 ;
        RECT 0.504 0.252 0.652 0.324 ;
        RECT 0.504 0.252 0.576 0.684 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.052 0.144 1.156 0.216 ;
      LAYER M1 ;
        RECT 1.044 0.144 1.156 0.216 ;
        RECT 0.072 0.756 0.92 0.828 ;
        RECT 0.052 0.144 0.252 0.216 ;
        RECT 0.072 0.144 0.144 0.828 ;
      LAYER V1 ;
        RECT 0.072 0.144 0.144 0.216 ;
        RECT 1.064 0.144 1.136 0.216 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.268 0.432 1.028 0.504 ;
      LAYER M1 ;
        RECT 0.936 0.412 1.008 0.596 ;
        RECT 0.288 0.412 0.36 0.596 ;
      LAYER V1 ;
        RECT 0.288 0.432 0.36 0.504 ;
        RECT 0.936 0.432 1.008 0.504 ;
    END
  END B1
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.568 0.972 ;
      RECT 0.376 0.108 0.92 0.18 ;
  END
END AOI32_xp67_75t

MACRO AOI331_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI331_xp33_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.136 0.576 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.136 0.36 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.668 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 0.804 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.016 0.756 1.572 0.828 ;
      RECT 0.368 0.9 1.356 0.972 ;
  END
END AOI331_xp33_75t

MACRO AOI332_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI332_xp33_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.136 0.576 0.656 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.136 0.36 0.656 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.668 0.756 2.088 0.828 ;
        RECT 2.016 0.108 2.088 0.828 ;
        RECT 0.804 0.108 2.088 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.016 0.9 2.008 0.972 ;
      RECT 0.368 0.756 1.356 0.828 ;
  END
END AOI332_xp33_75t

MACRO AOI333_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI333_xp33_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.28 2.088 0.656 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.656 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.656 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.136 0.576 0.656 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.136 0.36 0.656 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.652 0.756 2.304 0.828 ;
        RECT 2.232 0.108 2.304 0.828 ;
        RECT 0.804 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.016 0.9 2.06 0.972 ;
      RECT 0.376 0.756 1.36 0.828 ;
  END
END AOI333_xp33_75t

MACRO AOI33_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33_x1_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.748 1.084 0.82 ;
        RECT 0.936 0.404 1.084 0.476 ;
        RECT 0.936 0.404 1.008 0.82 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.508 0.748 1.656 0.82 ;
        RECT 1.584 0.404 1.656 0.82 ;
        RECT 1.508 0.404 1.656 0.476 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.088 0.604 2.304 0.676 ;
        RECT 2.232 0.404 2.304 0.676 ;
        RECT 2.088 0.604 2.16 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.26 2.52 0.656 ;
        RECT 2.372 0.26 2.52 0.332 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.664 0.28 2.736 0.656 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.32 0.756 2.952 0.828 ;
        RECT 2.88 0.108 2.952 0.828 ;
        RECT 1.672 0.108 2.952 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.592 0.9 2.648 0.972 ;
      RECT 1.024 0.252 2 0.324 ;
      RECT 0.376 0.108 1.352 0.18 ;
  END
END AOI33_x1_75t

MACRO AOI33_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33_xp33_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.136 0.36 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.136 0.576 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.656 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.656 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.656 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.756 1.656 0.828 ;
        RECT 1.584 0.108 1.656 0.828 ;
        RECT 0.804 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.9 1.352 0.972 ;
  END
END AOI33_xp33_75t

MACRO ASYNC_DFFH_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ASYNC_DFFH_x1_75t 0 0 ;
  SIZE 5.616 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.728 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.352 ;
        RECT 0.396 0.136 0.468 0.352 ;
        RECT 0.288 0.728 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.504 1.16 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.344 0.9 5.544 0.972 ;
        RECT 5.472 0.108 5.544 0.972 ;
        RECT 5.344 0.108 5.544 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.616 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.616 0.036 ;
    END
  END VSS
  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.528 0.432 4.268 0.504 ;
      LAYER M1 ;
        RECT 4.176 0.412 4.248 0.672 ;
        RECT 2.448 0.72 2.672 0.792 ;
        RECT 2.448 0.432 2.648 0.504 ;
        RECT 2.448 0.432 2.52 0.792 ;
      LAYER V1 ;
        RECT 2.548 0.432 2.62 0.504 ;
        RECT 4.176 0.432 4.248 0.504 ;
    END
  END RESET
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.132 0.288 4.268 0.36 ;
      LAYER M1 ;
        RECT 3.096 0.288 3.244 0.36 ;
        RECT 3.096 0.288 3.168 0.692 ;
      LAYER V1 ;
        RECT 3.152 0.288 3.224 0.36 ;
    END
  END SET
  OBS
    LAYER M1 ;
      RECT 3.852 0.864 4.032 0.936 ;
      RECT 3.852 0.144 3.924 0.936 ;
      RECT 3.672 0.12 3.744 0.868 ;
      RECT 3.432 0.12 3.744 0.192 ;
      RECT 2.232 0.864 3.08 0.936 ;
      RECT 2.772 0.232 2.844 0.936 ;
      RECT 2.232 0.656 2.304 0.936 ;
      RECT 1.672 0.9 2.016 0.972 ;
      RECT 1.944 0.288 2.016 0.972 ;
      RECT 1.944 0.288 2.188 0.36 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.072 0.9 0.272 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.072 0.576 0.188 0.648 ;
      RECT 0.072 0.108 0.272 0.18 ;
      RECT 5.256 0.36 5.328 0.668 ;
      RECT 4.68 0.144 4.808 0.216 ;
      RECT 4.392 0.412 4.464 0.672 ;
      RECT 3.528 0.388 3.6 0.812 ;
      RECT 3.316 0.396 3.388 0.668 ;
      RECT 3.112 0.144 3.276 0.216 ;
      RECT 2.916 0.268 2.988 0.532 ;
      RECT 1.66 0.108 2.432 0.18 ;
      RECT 1.8 0.476 1.872 0.668 ;
      RECT 1.584 0.48 1.656 0.812 ;
      RECT 1.476 0.216 1.548 0.404 ;
      RECT 1.368 0.48 1.44 0.668 ;
      RECT 0.568 0.424 0.64 0.668 ;
    LAYER M2 ;
      RECT 3.652 0.576 5.348 0.648 ;
      RECT 3.132 0.144 4.792 0.216 ;
      RECT 2.964 0.864 4.032 0.936 ;
      RECT 0.7 0.72 3.704 0.792 ;
      RECT 0.076 0.576 3.408 0.648 ;
      RECT 1.456 0.288 3.008 0.36 ;
    LAYER V1 ;
      RECT 5.256 0.576 5.328 0.648 ;
      RECT 4.7 0.144 4.772 0.216 ;
      RECT 4.392 0.576 4.464 0.648 ;
      RECT 3.94 0.864 4.012 0.936 ;
      RECT 3.672 0.576 3.744 0.648 ;
      RECT 3.528 0.72 3.6 0.792 ;
      RECT 3.316 0.576 3.388 0.648 ;
      RECT 3.152 0.144 3.224 0.216 ;
      RECT 2.984 0.864 3.056 0.936 ;
      RECT 2.916 0.288 2.988 0.36 ;
      RECT 2.048 0.288 2.12 0.36 ;
      RECT 1.8 0.576 1.872 0.648 ;
      RECT 1.584 0.72 1.656 0.792 ;
      RECT 1.476 0.288 1.548 0.36 ;
      RECT 1.368 0.576 1.44 0.648 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.568 0.576 0.64 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END ASYNC_DFFH_x1_75t

MACRO ASYNC_DFFH_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ASYNC_DFFH_x2_75t 0 0 ;
  SIZE 5.832 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.728 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.352 ;
        RECT 0.396 0.136 0.468 0.352 ;
        RECT 0.288 0.728 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.504 1.16 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.344 0.9 5.544 0.972 ;
        RECT 5.472 0.108 5.544 0.972 ;
        RECT 5.344 0.108 5.544 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.832 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.832 0.036 ;
    END
  END VSS
  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 2.528 0.432 4.268 0.504 ;
      LAYER M1 ;
        RECT 4.176 0.412 4.248 0.672 ;
        RECT 2.448 0.72 2.672 0.792 ;
        RECT 2.448 0.432 2.648 0.504 ;
        RECT 2.448 0.432 2.52 0.792 ;
      LAYER V1 ;
        RECT 2.548 0.432 2.62 0.504 ;
        RECT 4.176 0.432 4.248 0.504 ;
    END
  END RESET
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 3.132 0.288 4.268 0.36 ;
      LAYER M1 ;
        RECT 3.096 0.288 3.244 0.36 ;
        RECT 3.096 0.288 3.168 0.692 ;
      LAYER V1 ;
        RECT 3.152 0.288 3.224 0.36 ;
    END
  END SET
  OBS
    LAYER M1 ;
      RECT 3.852 0.864 4.032 0.936 ;
      RECT 3.852 0.144 3.924 0.936 ;
      RECT 3.672 0.12 3.744 0.868 ;
      RECT 3.432 0.12 3.744 0.192 ;
      RECT 2.232 0.864 3.08 0.936 ;
      RECT 2.772 0.232 2.844 0.936 ;
      RECT 2.232 0.656 2.304 0.936 ;
      RECT 1.672 0.9 2.016 0.972 ;
      RECT 1.944 0.288 2.016 0.972 ;
      RECT 1.944 0.288 2.188 0.36 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.072 0.9 0.272 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.072 0.576 0.188 0.648 ;
      RECT 0.072 0.108 0.272 0.18 ;
      RECT 5.256 0.36 5.328 0.668 ;
      RECT 4.68 0.144 4.808 0.216 ;
      RECT 4.392 0.412 4.464 0.672 ;
      RECT 3.528 0.388 3.6 0.812 ;
      RECT 3.316 0.396 3.388 0.668 ;
      RECT 3.112 0.144 3.276 0.216 ;
      RECT 2.916 0.268 2.988 0.532 ;
      RECT 1.66 0.108 2.432 0.18 ;
      RECT 1.8 0.476 1.872 0.668 ;
      RECT 1.584 0.48 1.656 0.812 ;
      RECT 1.476 0.216 1.548 0.404 ;
      RECT 1.368 0.48 1.44 0.668 ;
      RECT 0.568 0.424 0.64 0.668 ;
    LAYER M2 ;
      RECT 3.652 0.576 5.348 0.648 ;
      RECT 3.132 0.144 4.792 0.216 ;
      RECT 2.964 0.864 4.032 0.936 ;
      RECT 0.7 0.72 3.704 0.792 ;
      RECT 0.076 0.576 3.408 0.648 ;
      RECT 1.456 0.288 3.008 0.36 ;
    LAYER V1 ;
      RECT 5.256 0.576 5.328 0.648 ;
      RECT 4.7 0.144 4.772 0.216 ;
      RECT 4.392 0.576 4.464 0.648 ;
      RECT 3.94 0.864 4.012 0.936 ;
      RECT 3.672 0.576 3.744 0.648 ;
      RECT 3.528 0.72 3.6 0.792 ;
      RECT 3.316 0.576 3.388 0.648 ;
      RECT 3.152 0.144 3.224 0.216 ;
      RECT 2.984 0.864 3.056 0.936 ;
      RECT 2.916 0.288 2.988 0.36 ;
      RECT 2.048 0.288 2.12 0.36 ;
      RECT 1.8 0.576 1.872 0.648 ;
      RECT 1.584 0.72 1.656 0.792 ;
      RECT 1.476 0.288 1.548 0.36 ;
      RECT 1.368 0.576 1.44 0.648 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.568 0.576 0.64 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END ASYNC_DFFH_x2_75t

MACRO BUF_x10_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x10_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.9 2.952 0.972 ;
        RECT 2.88 0.108 2.952 0.972 ;
        RECT 0.796 0.108 2.952 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 2.756 0.576 ;
      RECT 0.364 0.108 0.576 0.18 ;
  END
END BUF_x10_75t

MACRO BUF_x12_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x12_75t 0 0 ;
  SIZE 3.456 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.456 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.9 3.384 0.972 ;
        RECT 3.312 0.108 3.384 0.972 ;
        RECT 0.796 0.108 3.384 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 3.2 0.576 ;
      RECT 0.376 0.108 0.576 0.18 ;
  END
END BUF_x12_75t

MACRO BUF_x12f_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x12f_75t 0 0 ;
  SIZE 3.888 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.316 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.888 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.888 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 3.816 0.972 ;
        RECT 3.744 0.108 3.816 0.972 ;
        RECT 1.24 0.108 3.816 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 1.116 0.972 ;
      RECT 1.044 0.108 1.116 0.972 ;
      RECT 1.044 0.504 1.244 0.576 ;
      RECT 0.376 0.108 1.116 0.18 ;
  END
END BUF_x12f_75t

MACRO BUF_x16f_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x16f_75t 0 0 ;
  SIZE 4.752 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.316 0.576 ;
        RECT 0.072 0.888 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.192 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.752 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.752 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 4.68 0.972 ;
        RECT 4.608 0.108 4.68 0.972 ;
        RECT 1.24 0.108 4.68 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.936 0.504 4.496 0.576 ;
      RECT 0.376 0.108 1.008 0.18 ;
  END
END BUF_x16f_75t

MACRO BUF_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x1_75t 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.58 0.108 0.792 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 0.596 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUF_x1_75t

MACRO BUF_x24_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x24_75t 0 0 ;
  SIZE 6.48 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 6.48 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.48 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 6.408 0.972 ;
        RECT 6.336 0.108 6.408 0.972 ;
        RECT 1.24 0.108 6.408 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.936 0.504 6.212 0.576 ;
      RECT 0.376 0.108 1.008 0.18 ;
  END
END BUF_x24_75t

MACRO BUF_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x2_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.58 0.108 1.008 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 0.812 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUF_x2_75t

MACRO BUF_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x3_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.58 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 1.04 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUF_x3_75t

MACRO BUF_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x4_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 1.428 0.972 ;
        RECT 1.356 0.108 1.428 0.972 ;
        RECT 0.58 0.108 1.428 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 1.256 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUF_x4_75t

MACRO BUF_x4f_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x4f_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.392 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.796 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.796 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 1.468 0.576 ;
      RECT 0.364 0.108 0.576 0.18 ;
  END
END BUF_x4f_75t

MACRO BUF_x5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x5_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.58 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 1.472 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUF_x5_75t

MACRO BUF_x6f_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x6f_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 2.088 0.972 ;
        RECT 2.016 0.108 2.088 0.972 ;
        RECT 0.808 0.108 2.088 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 1.892 0.576 ;
      RECT 0.376 0.108 0.576 0.18 ;
  END
END BUF_x6f_75t

MACRO BUF_x8_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_x8_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.392 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 2.52 0.972 ;
        RECT 2.448 0.108 2.52 0.972 ;
        RECT 0.808 0.108 2.52 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.364 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 2.324 0.576 ;
      RECT 0.364 0.108 0.576 0.18 ;
  END
END BUF_x8_75t

MACRO BUF_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_xp33_75t 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.58 0.108 0.792 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 0.596 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUF_xp33_75t

MACRO BUF_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_xp67_75t 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.292 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.58 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.58 0.108 0.792 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.48 0.972 ;
      RECT 0.408 0.108 0.48 0.972 ;
      RECT 0.408 0.504 0.596 0.576 ;
      RECT 0.16 0.108 0.48 0.18 ;
  END
END BUF_xp67_75t

MACRO DECAP_x10_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAP_x10_75t 0 0 ;
  SIZE 4.752 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.752 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.752 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.232 0.18 2.304 0.6 ;
      RECT 2.232 0.18 4.592 0.252 ;
      RECT 0.16 0.828 2.52 0.9 ;
      RECT 2.448 0.484 2.52 0.9 ;
  END
END DECAP_x10_75t

MACRO DECAP_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAP_x1_75t 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.376 0.828 0.576 0.9 ;
      RECT 0.504 0.484 0.576 0.9 ;
      RECT 0.288 0.18 0.36 0.6 ;
      RECT 0.288 0.18 0.488 0.252 ;
  END
END DECAP_x1_75t

MACRO DECAP_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAP_x2_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.504 0.18 0.576 0.6 ;
      RECT 0.504 0.18 1.136 0.252 ;
      RECT 0.16 0.828 0.792 0.9 ;
      RECT 0.72 0.484 0.792 0.9 ;
  END
END DECAP_x2_75t

MACRO DECAP_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAP_x4_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.936 0.18 1.008 0.6 ;
      RECT 0.936 0.18 2 0.252 ;
      RECT 0.16 0.828 1.224 0.9 ;
      RECT 1.152 0.484 1.224 0.9 ;
  END
END DECAP_x4_75t

MACRO DECAP_x6_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAP_x6_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.368 0.18 1.44 0.6 ;
      RECT 1.368 0.18 2.864 0.252 ;
      RECT 0.16 0.828 1.656 0.9 ;
      RECT 1.584 0.484 1.656 0.9 ;
  END
END DECAP_x6_75t

MACRO DFFHQN_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQN_x1_75t 0 0 ;
  SIZE 4.32 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.656 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.424 ;
        RECT 0.396 0.136 0.468 0.424 ;
        RECT 0.288 0.656 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.504 1.16 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.048 0.9 4.248 0.972 ;
        RECT 4.176 0.108 4.248 0.972 ;
        RECT 4.048 0.108 4.248 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.32 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.4 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.096 0.108 3.168 0.476 ;
      RECT 3.096 0.108 3.816 0.18 ;
      RECT 2.752 0.896 2.952 0.968 ;
      RECT 2.88 0.108 2.952 0.968 ;
      RECT 2.88 0.612 3.6 0.684 ;
      RECT 3.528 0.468 3.6 0.684 ;
      RECT 3.312 0.468 3.384 0.684 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 2.304 0.9 2.52 0.972 ;
      RECT 2.448 0.324 2.52 0.972 ;
      RECT 1.984 0.324 2.52 0.396 ;
      RECT 2.34 0.18 2.412 0.396 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.304 0.56 ;
      RECT 1.672 0.108 1.872 0.18 ;
      RECT 1.26 0.504 1.332 0.812 ;
      RECT 1.26 0.504 1.468 0.576 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.576 0.188 0.648 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.96 0.36 4.032 0.668 ;
      RECT 2.664 0.404 2.736 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.668 ;
      RECT 0.568 0.424 0.64 0.668 ;
    LAYER M2 ;
      RECT 3.508 0.576 4.052 0.648 ;
      RECT 0.076 0.576 2.756 0.648 ;
      RECT 0.7 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 3.96 0.576 4.032 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.664 0.576 2.736 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.26 0.72 1.332 0.792 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.568 0.576 0.64 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END DFFHQN_x1_75t

MACRO DFFHQN_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQN_x2_75t 0 0 ;
  SIZE 4.536 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.656 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.424 ;
        RECT 0.396 0.136 0.468 0.424 ;
        RECT 0.288 0.656 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.504 1.16 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.048 0.864 4.468 0.936 ;
        RECT 4.396 0.144 4.468 0.936 ;
        RECT 4.048 0.144 4.468 0.216 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.536 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.536 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.4 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.096 0.108 3.168 0.476 ;
      RECT 3.096 0.108 3.816 0.18 ;
      RECT 2.752 0.896 2.952 0.968 ;
      RECT 2.88 0.108 2.952 0.968 ;
      RECT 2.88 0.612 3.6 0.684 ;
      RECT 3.528 0.468 3.6 0.684 ;
      RECT 3.312 0.468 3.384 0.684 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 2.304 0.9 2.52 0.972 ;
      RECT 2.448 0.324 2.52 0.972 ;
      RECT 1.984 0.324 2.52 0.396 ;
      RECT 2.34 0.18 2.412 0.396 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.304 0.56 ;
      RECT 1.672 0.108 1.872 0.18 ;
      RECT 1.26 0.504 1.332 0.812 ;
      RECT 1.26 0.504 1.468 0.576 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.576 0.188 0.648 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.96 0.36 4.032 0.668 ;
      RECT 2.664 0.404 2.736 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.668 ;
      RECT 0.568 0.424 0.64 0.668 ;
    LAYER M2 ;
      RECT 3.508 0.576 4.052 0.648 ;
      RECT 0.076 0.576 2.756 0.648 ;
      RECT 0.7 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 3.96 0.576 4.032 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.664 0.576 2.736 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.26 0.72 1.332 0.792 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.568 0.576 0.64 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END DFFHQN_x2_75t

MACRO DFFHQN_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQN_x3_75t 0 0 ;
  SIZE 4.752 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.656 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.424 ;
        RECT 0.396 0.136 0.468 0.424 ;
        RECT 0.288 0.656 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.504 1.16 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.048 0.9 4.684 0.972 ;
        RECT 4.612 0.108 4.684 0.972 ;
        RECT 4.048 0.108 4.684 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.752 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.752 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.4 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.096 0.108 3.168 0.476 ;
      RECT 3.096 0.108 3.816 0.18 ;
      RECT 2.752 0.896 2.952 0.968 ;
      RECT 2.88 0.108 2.952 0.968 ;
      RECT 2.88 0.612 3.6 0.684 ;
      RECT 3.528 0.468 3.6 0.684 ;
      RECT 3.312 0.468 3.384 0.684 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 2.304 0.9 2.52 0.972 ;
      RECT 2.448 0.324 2.52 0.972 ;
      RECT 1.984 0.324 2.52 0.396 ;
      RECT 2.34 0.18 2.412 0.396 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.304 0.56 ;
      RECT 1.672 0.108 1.872 0.18 ;
      RECT 1.26 0.504 1.332 0.812 ;
      RECT 1.26 0.504 1.468 0.576 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.576 0.188 0.648 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.96 0.488 4.032 0.668 ;
      RECT 2.664 0.404 2.736 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.668 ;
      RECT 0.568 0.424 0.64 0.668 ;
    LAYER M2 ;
      RECT 3.508 0.576 4.052 0.648 ;
      RECT 0.076 0.576 2.756 0.648 ;
      RECT 0.7 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 3.96 0.576 4.032 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.664 0.576 2.736 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.26 0.72 1.332 0.792 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.568 0.576 0.64 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END DFFHQN_x3_75t

MACRO DFFHQ_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQ_x4_75t 0 0 ;
  SIZE 5.4 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.656 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.424 ;
        RECT 0.396 0.136 0.468 0.424 ;
        RECT 0.288 0.656 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.504 1.16 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5 0.9 5.332 0.972 ;
        RECT 5.252 0.108 5.332 0.972 ;
        RECT 4.5 0.108 5.332 0.18 ;
        RECT 4.5 0.804 4.572 0.972 ;
        RECT 4.5 0.108 4.572 0.276 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.4 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.4 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.048 0.9 4.392 0.972 ;
      RECT 4.32 0.108 4.392 0.972 ;
      RECT 4.32 0.508 4.7 0.58 ;
      RECT 4.048 0.108 4.392 0.18 ;
      RECT 3.4 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.096 0.108 3.168 0.476 ;
      RECT 3.096 0.108 3.816 0.18 ;
      RECT 2.752 0.896 2.952 0.968 ;
      RECT 2.88 0.108 2.952 0.968 ;
      RECT 2.88 0.612 3.6 0.684 ;
      RECT 3.528 0.468 3.6 0.684 ;
      RECT 3.312 0.468 3.384 0.684 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 2.304 0.9 2.52 0.972 ;
      RECT 2.448 0.324 2.52 0.972 ;
      RECT 1.984 0.324 2.52 0.396 ;
      RECT 2.34 0.18 2.412 0.396 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.324 0.56 ;
      RECT 1.672 0.108 1.872 0.18 ;
      RECT 1.26 0.504 1.332 0.812 ;
      RECT 1.26 0.504 1.468 0.576 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.576 0.188 0.648 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.96 0.488 4.032 0.668 ;
      RECT 2.664 0.404 2.736 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.668 ;
      RECT 0.568 0.424 0.64 0.668 ;
    LAYER M2 ;
      RECT 3.508 0.576 4.052 0.648 ;
      RECT 0.076 0.576 2.756 0.648 ;
      RECT 0.7 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 3.96 0.576 4.032 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.664 0.576 2.736 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.26 0.72 1.332 0.792 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.568 0.576 0.64 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END DFFHQ_x4_75t

MACRO DFFLQN_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQN_x1_75t 0 0 ;
  SIZE 4.32 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.656 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.424 ;
        RECT 0.396 0.136 0.468 0.424 ;
        RECT 0.288 0.656 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.9 1.3 0.972 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.048 0.9 4.248 0.972 ;
        RECT 4.176 0.108 4.248 0.972 ;
        RECT 4.048 0.108 4.248 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.32 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.4 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.096 0.108 3.168 0.476 ;
      RECT 3.096 0.108 3.816 0.18 ;
      RECT 2.752 0.9 2.952 0.972 ;
      RECT 2.88 0.108 2.952 0.972 ;
      RECT 2.88 0.612 3.6 0.684 ;
      RECT 3.528 0.468 3.6 0.684 ;
      RECT 3.312 0.468 3.384 0.684 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 2.304 0.9 2.52 0.972 ;
      RECT 2.448 0.324 2.52 0.972 ;
      RECT 1.984 0.324 2.52 0.396 ;
      RECT 2.34 0.136 2.412 0.396 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.324 0.56 ;
      RECT 1.672 0.108 1.872 0.18 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.58 0.72 0.792 0.792 ;
      RECT 0.72 0.504 0.792 0.792 ;
      RECT 0.484 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.96 0.36 4.032 0.668 ;
      RECT 2.664 0.396 2.736 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.668 ;
      RECT 1.368 0.504 1.44 0.812 ;
    LAYER M2 ;
      RECT 3.508 0.576 4.052 0.648 ;
      RECT 0.916 0.576 2.756 0.648 ;
      RECT 0.076 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 3.96 0.576 4.032 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.664 0.576 2.736 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.576 1.008 0.648 ;
      RECT 0.6 0.72 0.672 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END DFFLQN_x1_75t

MACRO DFFLQN_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQN_x2_75t 0 0 ;
  SIZE 4.536 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.656 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.424 ;
        RECT 0.396 0.136 0.468 0.424 ;
        RECT 0.288 0.656 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.9 1.3 0.972 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.048 0.9 4.46 0.972 ;
        RECT 4.388 0.108 4.46 0.972 ;
        RECT 4.048 0.108 4.46 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.536 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.536 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.4 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.096 0.108 3.168 0.476 ;
      RECT 3.096 0.108 3.816 0.18 ;
      RECT 2.752 0.9 2.952 0.972 ;
      RECT 2.88 0.108 2.952 0.972 ;
      RECT 2.88 0.612 3.6 0.684 ;
      RECT 3.528 0.468 3.6 0.684 ;
      RECT 3.312 0.468 3.384 0.684 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 2.304 0.9 2.52 0.972 ;
      RECT 2.448 0.324 2.52 0.972 ;
      RECT 1.984 0.324 2.52 0.396 ;
      RECT 2.34 0.136 2.412 0.396 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.324 0.56 ;
      RECT 1.672 0.108 1.872 0.18 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.58 0.72 0.792 0.792 ;
      RECT 0.72 0.504 0.792 0.792 ;
      RECT 0.484 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.96 0.36 4.032 0.668 ;
      RECT 2.664 0.396 2.736 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.668 ;
      RECT 1.368 0.504 1.44 0.812 ;
    LAYER M2 ;
      RECT 3.508 0.576 4.052 0.648 ;
      RECT 0.916 0.576 2.756 0.648 ;
      RECT 0.076 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 3.96 0.576 4.032 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.664 0.576 2.736 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.576 1.008 0.648 ;
      RECT 0.6 0.72 0.672 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END DFFLQN_x2_75t

MACRO DFFLQN_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQN_x3_75t 0 0 ;
  SIZE 4.752 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.656 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.424 ;
        RECT 0.396 0.136 0.468 0.424 ;
        RECT 0.288 0.656 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.9 1.3 0.972 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.048 0.9 4.684 0.972 ;
        RECT 4.612 0.108 4.684 0.972 ;
        RECT 4.044 0.108 4.684 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.752 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.752 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 3.4 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.096 0.108 3.168 0.476 ;
      RECT 3.096 0.108 3.816 0.18 ;
      RECT 2.752 0.9 2.952 0.972 ;
      RECT 2.88 0.108 2.952 0.972 ;
      RECT 2.88 0.612 3.6 0.684 ;
      RECT 3.528 0.468 3.6 0.684 ;
      RECT 3.312 0.468 3.384 0.684 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 2.304 0.9 2.52 0.972 ;
      RECT 2.448 0.324 2.52 0.972 ;
      RECT 1.984 0.324 2.52 0.396 ;
      RECT 2.34 0.136 2.412 0.396 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.324 0.56 ;
      RECT 1.672 0.108 1.872 0.18 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.58 0.72 0.792 0.792 ;
      RECT 0.72 0.504 0.792 0.792 ;
      RECT 0.484 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.96 0.36 4.032 0.668 ;
      RECT 2.664 0.396 2.736 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.668 ;
      RECT 1.368 0.504 1.44 0.812 ;
    LAYER M2 ;
      RECT 3.508 0.576 4.052 0.648 ;
      RECT 0.916 0.576 2.756 0.648 ;
      RECT 0.076 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 3.96 0.576 4.032 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.664 0.576 2.736 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.576 1.008 0.648 ;
      RECT 0.6 0.72 0.672 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END DFFLQN_x3_75t

MACRO DFFLQ_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFLQ_x4_75t 0 0 ;
  SIZE 5.4 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.656 0.468 0.944 ;
        RECT 0.288 0.28 0.468 0.424 ;
        RECT 0.396 0.136 0.468 0.424 ;
        RECT 0.288 0.656 0.468 0.8 ;
        RECT 0.288 0.28 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.9 1.3 0.972 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.972 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 4.5 0.9 5.332 0.972 ;
        RECT 5.252 0.108 5.332 0.972 ;
        RECT 4.5 0.108 5.332 0.18 ;
        RECT 4.5 0.804 4.572 0.972 ;
        RECT 4.5 0.108 4.572 0.276 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.4 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.4 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.048 0.9 4.392 0.972 ;
      RECT 4.32 0.108 4.392 0.972 ;
      RECT 4.32 0.508 4.7 0.58 ;
      RECT 4.048 0.108 4.392 0.18 ;
      RECT 3.4 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.096 0.108 3.168 0.476 ;
      RECT 3.096 0.108 3.816 0.18 ;
      RECT 2.752 0.9 2.952 0.972 ;
      RECT 2.88 0.108 2.952 0.972 ;
      RECT 2.88 0.612 3.6 0.684 ;
      RECT 3.528 0.468 3.6 0.684 ;
      RECT 3.312 0.468 3.384 0.684 ;
      RECT 2.536 0.108 2.952 0.18 ;
      RECT 2.304 0.9 2.52 0.972 ;
      RECT 2.448 0.324 2.52 0.972 ;
      RECT 1.984 0.324 2.52 0.396 ;
      RECT 2.34 0.136 2.412 0.396 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.324 0.56 ;
      RECT 1.672 0.108 1.872 0.18 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.58 0.72 0.792 0.792 ;
      RECT 0.72 0.504 0.792 0.792 ;
      RECT 0.484 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.96 0.488 4.032 0.668 ;
      RECT 2.664 0.396 2.736 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.668 ;
      RECT 1.368 0.504 1.44 0.812 ;
    LAYER M2 ;
      RECT 3.508 0.576 4.052 0.648 ;
      RECT 0.916 0.576 2.756 0.648 ;
      RECT 0.076 0.72 2.108 0.792 ;
    LAYER V1 ;
      RECT 3.96 0.576 4.032 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.664 0.576 2.736 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.576 1.008 0.648 ;
      RECT 0.6 0.72 0.672 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END DFFLQ_x4_75t

MACRO DHL_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHL_x1_75t 0 0 ;
  SIZE 3.24 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.612 0.468 0.944 ;
        RECT 0.288 0.324 0.468 0.468 ;
        RECT 0.396 0.136 0.468 0.468 ;
        RECT 0.288 0.612 0.468 0.756 ;
        RECT 0.288 0.324 0.36 0.756 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.944 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.968 0.9 3.168 0.972 ;
        RECT 3.096 0.108 3.168 0.972 ;
        RECT 2.968 0.108 3.168 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.24 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.32 0.9 2.52 0.972 ;
      RECT 2.448 0.108 2.52 0.972 ;
      RECT 2.016 0.108 2.088 0.384 ;
      RECT 2.016 0.108 2.52 0.18 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.484 2.324 0.556 ;
      RECT 1.656 0.108 1.872 0.18 ;
      RECT 1.368 0.756 1.516 0.828 ;
      RECT 1.368 0.424 1.44 0.828 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.592 0.72 0.792 0.792 ;
      RECT 0.72 0.504 0.792 0.792 ;
      RECT 0.552 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 2.88 0.488 2.952 0.668 ;
      RECT 2.016 0.656 2.088 0.828 ;
      RECT 1.584 0.424 1.656 0.684 ;
    LAYER M2 ;
      RECT 1.8 0.576 2.972 0.648 ;
      RECT 0.076 0.72 2.108 0.792 ;
      RECT 0.916 0.576 1.656 0.648 ;
    LAYER V1 ;
      RECT 2.88 0.576 2.952 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.8 0.576 1.872 0.648 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.576 1.008 0.648 ;
      RECT 0.612 0.72 0.684 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END DHL_x1_75t

MACRO DHL_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHL_x2_75t 0 0 ;
  SIZE 3.456 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.612 0.468 0.944 ;
        RECT 0.288 0.324 0.468 0.468 ;
        RECT 0.396 0.136 0.468 0.468 ;
        RECT 0.288 0.612 0.468 0.756 ;
        RECT 0.288 0.324 0.36 0.756 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.944 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.964 0.864 3.4 0.936 ;
        RECT 3.328 0.144 3.4 0.936 ;
        RECT 2.968 0.144 3.4 0.216 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.456 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.32 0.9 2.52 0.972 ;
      RECT 2.448 0.108 2.52 0.972 ;
      RECT 2.016 0.108 2.088 0.384 ;
      RECT 2.016 0.108 2.52 0.18 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.484 2.324 0.556 ;
      RECT 1.656 0.108 1.872 0.18 ;
      RECT 1.368 0.756 1.516 0.828 ;
      RECT 1.368 0.424 1.44 0.828 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.592 0.72 0.792 0.792 ;
      RECT 0.72 0.504 0.792 0.792 ;
      RECT 0.552 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.096 0.36 3.168 0.668 ;
      RECT 2.88 0.36 2.952 0.668 ;
      RECT 2.016 0.656 2.088 0.828 ;
      RECT 1.584 0.424 1.656 0.684 ;
    LAYER M2 ;
      RECT 1.8 0.576 3.188 0.648 ;
      RECT 0.076 0.72 2.108 0.792 ;
      RECT 0.916 0.576 1.656 0.648 ;
    LAYER V1 ;
      RECT 3.096 0.576 3.168 0.648 ;
      RECT 2.88 0.576 2.952 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.8 0.576 1.872 0.648 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.576 1.008 0.648 ;
      RECT 0.612 0.72 0.684 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END DHL_x2_75t

MACRO DHL_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHL_x3_75t 0 0 ;
  SIZE 3.672 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.612 0.468 0.944 ;
        RECT 0.288 0.324 0.468 0.468 ;
        RECT 0.396 0.136 0.468 0.468 ;
        RECT 0.288 0.612 0.468 0.756 ;
        RECT 0.288 0.324 0.36 0.756 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.944 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.752 0.9 3.6 0.972 ;
        RECT 3.528 0.108 3.6 0.972 ;
        RECT 2.752 0.108 3.6 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.672 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.672 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.32 0.9 2.52 0.972 ;
      RECT 2.448 0.108 2.52 0.972 ;
      RECT 2.016 0.108 2.088 0.384 ;
      RECT 2.016 0.108 2.52 0.18 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.484 2.324 0.556 ;
      RECT 1.656 0.108 1.872 0.18 ;
      RECT 1.368 0.756 1.516 0.828 ;
      RECT 1.368 0.424 1.44 0.828 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.592 0.72 0.792 0.792 ;
      RECT 0.72 0.504 0.792 0.792 ;
      RECT 0.552 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.312 0.36 3.384 0.668 ;
      RECT 3.096 0.36 3.168 0.668 ;
      RECT 2.88 0.36 2.952 0.668 ;
      RECT 2.016 0.656 2.088 0.828 ;
      RECT 1.584 0.424 1.656 0.684 ;
    LAYER M2 ;
      RECT 1.8 0.576 3.404 0.648 ;
      RECT 0.076 0.72 2.108 0.792 ;
      RECT 0.916 0.576 1.656 0.648 ;
    LAYER V1 ;
      RECT 3.312 0.576 3.384 0.648 ;
      RECT 3.096 0.576 3.168 0.648 ;
      RECT 2.88 0.576 2.952 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.8 0.576 1.872 0.648 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.576 1.008 0.648 ;
      RECT 0.612 0.72 0.684 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END DHL_x3_75t

MACRO DLL_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLL_x1_75t 0 0 ;
  SIZE 3.24 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.612 0.468 0.944 ;
        RECT 0.288 0.324 0.468 0.468 ;
        RECT 0.396 0.136 0.468 0.468 ;
        RECT 0.288 0.612 0.468 0.756 ;
        RECT 0.288 0.324 0.36 0.756 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.9 1.3 0.972 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.972 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.968 0.9 3.168 0.972 ;
        RECT 3.096 0.108 3.168 0.972 ;
        RECT 2.94 0.108 3.168 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.24 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.32 0.9 2.52 0.972 ;
      RECT 2.448 0.108 2.52 0.972 ;
      RECT 2.016 0.108 2.088 0.388 ;
      RECT 2.016 0.108 2.52 0.18 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.32 0.56 ;
      RECT 1.656 0.108 1.872 0.18 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.592 0.756 0.792 0.828 ;
      RECT 0.72 0.504 0.792 0.828 ;
      RECT 0.552 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.576 0.188 0.648 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 2.88 0.424 2.952 0.8 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.8 ;
      RECT 1.368 0.424 1.44 0.812 ;
    LAYER M2 ;
      RECT 1.8 0.576 2.972 0.648 ;
      RECT 0.916 0.72 2.108 0.792 ;
      RECT 0.076 0.576 1.656 0.648 ;
    LAYER V1 ;
      RECT 2.88 0.576 2.952 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.8 0.576 1.872 0.648 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.72 1.008 0.792 ;
      RECT 0.72 0.576 0.792 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END DLL_x1_75t

MACRO DLL_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLL_x2_75t 0 0 ;
  SIZE 3.456 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.612 0.468 0.944 ;
        RECT 0.288 0.324 0.468 0.468 ;
        RECT 0.396 0.136 0.468 0.468 ;
        RECT 0.288 0.612 0.468 0.756 ;
        RECT 0.288 0.324 0.36 0.756 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.9 1.3 0.972 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.972 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.752 0.9 3.388 0.972 ;
        RECT 3.316 0.108 3.388 0.972 ;
        RECT 2.752 0.108 3.388 0.18 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.456 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.32 0.9 2.52 0.972 ;
      RECT 2.448 0.108 2.52 0.972 ;
      RECT 2.016 0.108 2.088 0.388 ;
      RECT 2.016 0.108 2.52 0.18 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.32 0.56 ;
      RECT 1.656 0.108 1.872 0.18 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.592 0.756 0.792 0.828 ;
      RECT 0.72 0.504 0.792 0.828 ;
      RECT 0.552 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.576 0.188 0.648 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.096 0.36 3.168 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.8 ;
      RECT 1.368 0.424 1.44 0.812 ;
    LAYER M2 ;
      RECT 1.8 0.576 3.2 0.648 ;
      RECT 0.916 0.72 2.108 0.792 ;
      RECT 0.076 0.576 1.656 0.648 ;
    LAYER V1 ;
      RECT 3.096 0.576 3.168 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.8 0.576 1.872 0.648 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.72 1.008 0.792 ;
      RECT 0.72 0.576 0.792 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END DLL_x2_75t

MACRO DLL_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLL_x3_75t 0 0 ;
  SIZE 3.672 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.612 0.468 0.944 ;
        RECT 0.288 0.324 0.468 0.468 ;
        RECT 0.396 0.136 0.468 0.468 ;
        RECT 0.288 0.612 0.468 0.756 ;
        RECT 0.288 0.324 0.36 0.756 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.9 1.3 0.972 ;
        RECT 1.152 0.108 1.3 0.18 ;
        RECT 1.152 0.108 1.224 0.972 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.968 0.864 3.604 0.936 ;
        RECT 3.528 0.144 3.604 0.936 ;
        RECT 2.968 0.144 3.604 0.216 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.672 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.672 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 2.32 0.9 2.52 0.972 ;
      RECT 2.448 0.108 2.52 0.972 ;
      RECT 2.016 0.108 2.088 0.388 ;
      RECT 2.016 0.108 2.52 0.18 ;
      RECT 1.456 0.9 1.872 0.972 ;
      RECT 1.8 0.108 1.872 0.972 ;
      RECT 1.8 0.488 2.32 0.56 ;
      RECT 1.656 0.108 1.872 0.18 ;
      RECT 0.592 0.9 1.008 0.972 ;
      RECT 0.936 0.108 1.008 0.972 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 0.592 0.756 0.792 0.828 ;
      RECT 0.72 0.504 0.792 0.828 ;
      RECT 0.552 0.504 0.792 0.576 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.576 0.188 0.648 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 3.096 0.36 3.168 0.668 ;
      RECT 2.016 0.66 2.088 0.812 ;
      RECT 1.584 0.424 1.656 0.8 ;
      RECT 1.368 0.424 1.44 0.812 ;
    LAYER M2 ;
      RECT 1.8 0.576 3.2 0.648 ;
      RECT 0.916 0.72 2.108 0.792 ;
      RECT 0.076 0.576 1.656 0.648 ;
    LAYER V1 ;
      RECT 3.096 0.576 3.168 0.648 ;
      RECT 2.016 0.72 2.088 0.792 ;
      RECT 1.8 0.576 1.872 0.648 ;
      RECT 1.584 0.576 1.656 0.648 ;
      RECT 1.368 0.72 1.44 0.792 ;
      RECT 0.936 0.72 1.008 0.792 ;
      RECT 0.72 0.576 0.792 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END DLL_x3_75t

MACRO FA_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA_x1_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.296 0.9 1.98 0.972 ;
        RECT 1.908 0.736 1.98 0.972 ;
        RECT 1.908 0.108 1.98 0.272 ;
        RECT 1.296 0.108 1.98 0.18 ;
        RECT 1.296 0.108 1.368 0.972 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.236 0.72 2.508 0.792 ;
      LAYER M1 ;
        RECT 2.396 0.72 2.52 0.792 ;
        RECT 2.448 0.484 2.52 0.792 ;
        RECT 1.532 0.72 1.656 0.792 ;
        RECT 1.584 0.484 1.656 0.792 ;
        RECT 0.236 0.72 0.36 0.792 ;
        RECT 0.288 0.484 0.36 0.792 ;
      LAYER V1 ;
        RECT 0.256 0.72 0.328 0.792 ;
        RECT 1.552 0.72 1.624 0.792 ;
        RECT 2.416 0.72 2.488 0.792 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.668 0.576 2.756 0.648 ;
      LAYER M1 ;
        RECT 2.664 0.484 2.736 0.668 ;
        RECT 1.152 0.484 1.224 0.668 ;
        RECT 0.668 0.576 0.792 0.648 ;
        RECT 0.72 0.484 0.792 0.648 ;
      LAYER V1 ;
        RECT 0.688 0.576 0.76 0.648 ;
        RECT 1.152 0.576 1.224 0.648 ;
        RECT 2.664 0.576 2.736 0.648 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.916 0.432 2.348 0.504 ;
      LAYER M1 ;
        RECT 2.232 0.432 2.348 0.504 ;
        RECT 2.232 0.432 2.304 0.596 ;
        RECT 1.8 0.412 1.872 0.596 ;
        RECT 0.904 0.432 1.052 0.504 ;
        RECT 0.936 0.432 1.008 0.596 ;
      LAYER V1 ;
        RECT 0.936 0.432 1.008 0.504 ;
        RECT 1.8 0.432 1.872 0.504 ;
        RECT 2.256 0.432 2.328 0.504 ;
    END
  END CI
  PIN CON
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.512 0.288 2.172 0.36 ;
      LAYER M1 ;
        RECT 2.06 0.288 2.172 0.36 ;
        RECT 2.016 0.36 2.132 0.432 ;
        RECT 2.016 0.36 2.088 0.596 ;
        RECT 0.496 0.288 1.128 0.36 ;
        RECT 0.496 0.756 0.92 0.828 ;
        RECT 0.496 0.288 0.568 0.828 ;
      LAYER V1 ;
        RECT 0.532 0.288 0.604 0.36 ;
        RECT 2.08 0.288 2.152 0.36 ;
    END
  END CON
  OBS
    LAYER M1 ;
      RECT 2.104 0.108 2.648 0.18 ;
      RECT 2.104 0.9 2.648 0.972 ;
      RECT 0.16 0.108 1.136 0.18 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END FA_x1_75t

MACRO FILLER_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER_75t 0 0 ;
  SIZE 0.432 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.432 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.432 0.036 ;
    END
  END VSS
END FILLER_75t

MACRO FILLER_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER_xp5_75t 0 0 ;
  SIZE 0.216 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.216 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.216 0.036 ;
    END
  END VSS
END FILLER_xp5_75t

MACRO HA_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HA_x1_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.432 2.252 0.504 ;
        RECT 2.016 0.432 2.088 0.704 ;
        RECT 1.368 0.412 1.44 0.596 ;
        RECT 0.72 0.412 0.792 0.596 ;
      LAYER M2 ;
        RECT 0.7 0.432 2.252 0.504 ;
      LAYER V1 ;
        RECT 0.72 0.432 0.792 0.504 ;
        RECT 1.368 0.432 1.44 0.504 ;
        RECT 2.16 0.432 2.232 0.504 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.288 1.964 0.36 ;
        RECT 1.8 0.288 1.872 0.668 ;
        RECT 0.936 0.288 1.136 0.36 ;
        RECT 0.936 0.288 1.008 0.596 ;
      LAYER M2 ;
        RECT 1.024 0.288 1.964 0.36 ;
      LAYER V1 ;
        RECT 1.044 0.288 1.116 0.36 ;
        RECT 1.872 0.288 1.944 0.36 ;
    END
  END B
  PIN CON
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.512 0.9 2.304 0.972 ;
        RECT 1.512 0.556 1.584 0.972 ;
        RECT 1.656 0.34 1.728 0.668 ;
        RECT 0.224 0.392 0.296 0.668 ;
      LAYER M2 ;
        RECT 0.204 0.576 2.324 0.648 ;
      LAYER V1 ;
        RECT 0.224 0.576 0.296 0.648 ;
        RECT 1.512 0.576 1.584 0.648 ;
        RECT 1.656 0.576 1.728 0.648 ;
    END
  END CON
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.864 1.172 0.936 ;
        RECT 0.352 0.864 0.516 0.936 ;
        RECT 0.444 0.34 0.516 0.936 ;
      LAYER M2 ;
        RECT 0.352 0.864 1.172 0.936 ;
      LAYER V1 ;
        RECT 0.372 0.864 0.444 0.936 ;
        RECT 1.044 0.864 1.116 0.936 ;
    END
  END SN
  OBS
    LAYER M1 ;
      RECT 2.284 0.144 2.432 0.216 ;
      RECT 1.456 0.108 2 0.18 ;
      RECT 0.808 0.72 1.4 0.792 ;
      RECT 1.024 0.144 1.172 0.216 ;
      RECT 0.592 0.144 0.74 0.216 ;
      RECT 0.16 0.144 0.308 0.216 ;
    LAYER M2 ;
      RECT 0.16 0.144 2.432 0.216 ;
    LAYER V1 ;
      RECT 2.34 0.144 2.412 0.216 ;
      RECT 1.044 0.144 1.116 0.216 ;
      RECT 0.612 0.144 0.684 0.216 ;
      RECT 0.18 0.144 0.252 0.216 ;
  END
END HA_x1_75t

MACRO HA_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HA_xp5_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.252 1.44 0.6 ;
        RECT 0.828 0.252 1.44 0.324 ;
        RECT 0.828 0.108 0.9 0.324 ;
        RECT 0.072 0.108 0.9 0.18 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.896 0.22 0.968 ;
        RECT 0.072 0.108 0.144 0.968 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.424 0.252 0.576 0.324 ;
    END
  END B
  PIN CON
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.756 1.656 0.828 ;
        RECT 1.584 0.484 1.656 0.828 ;
        RECT 0.376 0.9 0.72 0.972 ;
        RECT 0.648 0.3 0.72 0.972 ;
    END
  END CON
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.692 0.108 1.872 0.18 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 1.024 0.108 1.548 0.18 ;
  END
END HA_xp5_75t

MACRO HB1_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB1_xp67_75t 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.896 0.792 0.968 ;
        RECT 0.72 0.104 0.792 0.968 ;
        RECT 0.592 0.104 0.792 0.176 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.468 0.972 ;
      RECT 0.396 0.612 0.468 0.972 ;
      RECT 0.396 0.612 0.576 0.684 ;
      RECT 0.504 0.396 0.576 0.684 ;
      RECT 0.396 0.396 0.576 0.468 ;
      RECT 0.396 0.108 0.468 0.468 ;
      RECT 0.16 0.108 0.468 0.18 ;
  END
END HB1_xp67_75t

MACRO HB2_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB2_xp67_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.808 0.108 1.008 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.576 0.972 ;
      RECT 0.504 0.108 0.576 0.972 ;
      RECT 0.504 0.504 0.812 0.576 ;
      RECT 0.16 0.108 0.576 0.18 ;
  END
END HB2_xp67_75t

MACRO HB3_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB3_xp67_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 1.024 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.72 0.504 1.028 0.576 ;
      RECT 0.16 0.108 0.792 0.18 ;
  END
END HB3_xp67_75t

MACRO HB4_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HB4_xp67_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.324 0.22 0.396 ;
        RECT 0.072 0.324 0.144 0.828 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.24 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.72 0.504 1.244 0.576 ;
      RECT 0.16 0.108 0.792 0.18 ;
  END
END HB4_xp67_75t

MACRO ICG_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICG_x1_75t 0 0 ;
  SIZE 3.888 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.796 ;
    END
  END ENA
  PIN GCLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 3.596 0.9 3.816 0.972 ;
        RECT 3.744 0.108 3.816 0.972 ;
        RECT 3.516 0.108 3.816 0.18 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.796 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.888 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.888 0.036 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.916 0.576 2.54 0.648 ;
      LAYER M1 ;
        RECT 2.448 0.712 3.06 0.784 ;
        RECT 2.988 0.568 3.06 0.784 ;
        RECT 2.448 0.464 2.52 0.784 ;
        RECT 1.584 0.576 1.788 0.648 ;
        RECT 1.584 0.48 1.656 0.648 ;
        RECT 0.936 0.476 1.008 0.736 ;
      LAYER V1 ;
        RECT 0.936 0.576 1.008 0.648 ;
        RECT 1.656 0.576 1.728 0.648 ;
        RECT 2.448 0.576 2.52 0.648 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 2.752 0.888 3.384 0.96 ;
      RECT 3.312 0.752 3.384 0.96 ;
      RECT 3.312 0.752 3.6 0.824 ;
      RECT 3.528 0.252 3.6 0.824 ;
      RECT 2.968 0.252 3.6 0.324 ;
      RECT 1.024 0.892 1.468 0.964 ;
      RECT 1.396 0.108 1.468 0.964 ;
      RECT 1.396 0.724 1.892 0.796 ;
      RECT 3.312 0.396 3.384 0.588 ;
      RECT 2.664 0.108 2.736 0.588 ;
      RECT 2.664 0.396 3.384 0.468 ;
      RECT 1.24 0.108 2.736 0.18 ;
      RECT 2.236 0.892 2.436 0.964 ;
      RECT 2.236 0.308 2.308 0.964 ;
      RECT 2.236 0.308 2.436 0.38 ;
      RECT 1.872 0.896 2.088 0.968 ;
      RECT 2.012 0.292 2.088 0.968 ;
      RECT 1.568 0.292 2.088 0.364 ;
      RECT 1.152 0.72 1.296 0.792 ;
      RECT 1.152 0.288 1.224 0.792 ;
      RECT 0.148 0.896 0.792 0.968 ;
      RECT 0.72 0.108 0.792 0.968 ;
      RECT 0.356 0.108 0.792 0.18 ;
    LAYER M2 ;
      RECT 1.184 0.72 2.328 0.792 ;
    LAYER V1 ;
      RECT 2.236 0.72 2.308 0.792 ;
      RECT 1.204 0.72 1.276 0.792 ;
  END
END ICG_x1_75t

MACRO ICG_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICG_x2_75t 0 0 ;
  SIZE 4.104 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.796 ;
    END
  END ENA
  PIN GCLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 3.596 0.9 4.032 0.972 ;
        RECT 3.96 0.108 4.032 0.972 ;
        RECT 3.516 0.108 4.032 0.18 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.796 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.104 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.104 0.036 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.916 0.576 2.54 0.648 ;
      LAYER M1 ;
        RECT 2.448 0.712 3.06 0.784 ;
        RECT 2.988 0.568 3.06 0.784 ;
        RECT 2.448 0.464 2.52 0.784 ;
        RECT 1.584 0.576 1.788 0.648 ;
        RECT 1.584 0.48 1.656 0.648 ;
        RECT 0.936 0.476 1.008 0.736 ;
      LAYER V1 ;
        RECT 0.936 0.576 1.008 0.648 ;
        RECT 1.656 0.576 1.728 0.648 ;
        RECT 2.448 0.576 2.52 0.648 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 2.752 0.888 3.384 0.96 ;
      RECT 3.312 0.752 3.384 0.96 ;
      RECT 3.312 0.752 3.6 0.824 ;
      RECT 3.528 0.252 3.6 0.824 ;
      RECT 2.968 0.252 3.6 0.324 ;
      RECT 1.024 0.892 1.468 0.964 ;
      RECT 1.396 0.108 1.468 0.964 ;
      RECT 1.396 0.724 1.892 0.796 ;
      RECT 3.312 0.396 3.384 0.588 ;
      RECT 2.664 0.108 2.736 0.588 ;
      RECT 2.664 0.396 3.384 0.468 ;
      RECT 1.24 0.108 2.736 0.18 ;
      RECT 2.236 0.892 2.436 0.964 ;
      RECT 2.236 0.308 2.308 0.964 ;
      RECT 2.236 0.308 2.436 0.38 ;
      RECT 1.872 0.896 2.088 0.968 ;
      RECT 2.012 0.292 2.088 0.968 ;
      RECT 1.568 0.292 2.088 0.364 ;
      RECT 1.152 0.72 1.296 0.792 ;
      RECT 1.152 0.288 1.224 0.792 ;
      RECT 1.028 0.288 1.224 0.36 ;
      RECT 0.148 0.896 0.792 0.968 ;
      RECT 0.72 0.108 0.792 0.968 ;
      RECT 0.356 0.108 0.792 0.18 ;
    LAYER M2 ;
      RECT 1.184 0.72 2.328 0.792 ;
    LAYER V1 ;
      RECT 2.236 0.72 2.308 0.792 ;
      RECT 1.204 0.72 1.276 0.792 ;
  END
END ICG_x2_75t

MACRO ICG_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ICG_x3_75t 0 0 ;
  SIZE 4.32 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN ENA
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.28 0.36 0.796 ;
    END
  END ENA
  PIN GCLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 3.596 0.9 4.248 0.972 ;
        RECT 4.176 0.108 4.248 0.972 ;
        RECT 3.516 0.108 4.248 0.18 ;
    END
  END GCLK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.796 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.32 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
    END
  END VSS
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M2 ;
        RECT 0.916 0.576 2.54 0.648 ;
      LAYER M1 ;
        RECT 2.448 0.712 3.06 0.784 ;
        RECT 2.988 0.568 3.06 0.784 ;
        RECT 2.448 0.464 2.52 0.784 ;
        RECT 1.584 0.576 1.788 0.648 ;
        RECT 1.584 0.48 1.656 0.648 ;
        RECT 0.936 0.476 1.008 0.736 ;
      LAYER V1 ;
        RECT 0.936 0.576 1.008 0.648 ;
        RECT 1.656 0.576 1.728 0.648 ;
        RECT 2.448 0.576 2.52 0.648 ;
    END
  END CLK
  OBS
    LAYER M1 ;
      RECT 2.752 0.888 3.384 0.96 ;
      RECT 3.312 0.752 3.384 0.96 ;
      RECT 3.312 0.752 3.6 0.824 ;
      RECT 3.528 0.252 3.6 0.824 ;
      RECT 2.968 0.252 3.6 0.324 ;
      RECT 1.024 0.892 1.468 0.964 ;
      RECT 1.396 0.108 1.468 0.964 ;
      RECT 1.396 0.724 1.892 0.796 ;
      RECT 3.312 0.396 3.384 0.588 ;
      RECT 2.664 0.108 2.736 0.588 ;
      RECT 2.664 0.396 3.384 0.468 ;
      RECT 1.24 0.108 2.736 0.18 ;
      RECT 2.236 0.892 2.436 0.964 ;
      RECT 2.236 0.308 2.308 0.964 ;
      RECT 2.236 0.308 2.436 0.38 ;
      RECT 1.872 0.896 2.088 0.968 ;
      RECT 2.012 0.292 2.088 0.968 ;
      RECT 1.568 0.292 2.088 0.364 ;
      RECT 1.152 0.72 1.296 0.792 ;
      RECT 1.152 0.288 1.224 0.792 ;
      RECT 1.028 0.288 1.224 0.36 ;
      RECT 0.148 0.896 0.792 0.968 ;
      RECT 0.72 0.108 0.792 0.968 ;
      RECT 0.356 0.108 0.792 0.18 ;
    LAYER M2 ;
      RECT 1.184 0.72 2.328 0.792 ;
    LAYER V1 ;
      RECT 2.236 0.72 2.308 0.792 ;
      RECT 1.204 0.72 1.276 0.792 ;
  END
END ICG_x3_75t

MACRO INV_x11_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_x11_75t 0 0 ;
  SIZE 2.808 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.808 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 2.736 0.972 ;
        RECT 2.664 0.108 2.736 0.972 ;
        RECT 0.376 0.108 2.736 0.18 ;
    END
  END Y
END INV_x11_75t

MACRO INV_x13_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_x13_75t 0 0 ;
  SIZE 3.24 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.24 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 3.168 0.972 ;
        RECT 3.096 0.108 3.168 0.972 ;
        RECT 0.376 0.108 3.168 0.18 ;
    END
  END Y
END INV_x13_75t

MACRO INV_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_x1_75t 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.576 0.972 ;
        RECT 0.504 0.108 0.576 0.972 ;
        RECT 0.376 0.108 0.576 0.18 ;
    END
  END Y
END INV_x1_75t

MACRO INV_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_x2_75t 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.376 0.108 0.792 0.18 ;
    END
  END Y
END INV_x2_75t

MACRO INV_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_x3_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.008 0.972 ;
        RECT 0.936 0.108 1.008 0.972 ;
        RECT 0.376 0.108 1.008 0.18 ;
    END
  END Y
END INV_x3_75t

MACRO INV_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_x4_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.376 0.108 1.224 0.18 ;
    END
  END Y
END INV_x4_75t

MACRO INV_x5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_x5_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 0.376 0.108 1.44 0.18 ;
    END
  END Y
END INV_x5_75t

MACRO INV_x6_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_x6_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.376 0.108 1.656 0.18 ;
    END
  END Y
END INV_x6_75t

MACRO INV_x8_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_x8_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 2.088 0.972 ;
        RECT 2.016 0.108 2.088 0.972 ;
        RECT 0.376 0.108 2.088 0.18 ;
    END
  END Y
END INV_x8_75t

MACRO INV_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_xp33_75t 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.9 0.576 0.972 ;
        RECT 0.504 0.108 0.576 0.972 ;
        RECT 0.336 0.504 0.576 0.576 ;
        RECT 0.428 0.108 0.576 0.18 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
END INV_xp33_75t

MACRO INV_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_xp67_75t 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.9 0.576 0.972 ;
        RECT 0.504 0.108 0.576 0.972 ;
        RECT 0.336 0.504 0.576 0.576 ;
        RECT 0.428 0.108 0.576 0.18 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
END INV_xp67_75t

MACRO MAJI_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJI_xp5_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.224 0.424 1.296 0.656 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.504 1.028 0.576 ;
        RECT 0.072 0.756 0.792 0.828 ;
        RECT 0.72 0.504 0.792 0.828 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.136 0.144 0.828 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.26 0.652 0.332 ;
        RECT 0.504 0.26 0.576 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.02 0.756 1.444 0.828 ;
        RECT 1.372 0.252 1.444 0.828 ;
        RECT 1.02 0.252 1.444 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.108 1.352 0.18 ;
      RECT 0.376 0.9 1.352 0.972 ;
  END
END MAJI_xp5_75t

MACRO MAJ_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJ_x2_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.424 0.288 0.656 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.756 1.332 0.828 ;
        RECT 1.26 0.424 1.332 0.828 ;
        RECT 1.132 0.504 1.332 0.576 ;
        RECT 0.592 0.504 0.664 0.828 ;
        RECT 0.484 0.504 0.664 0.576 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.764 0.612 1.008 0.684 ;
        RECT 0.936 0.396 1.008 0.684 ;
        RECT 0.764 0.396 1.008 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.456 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.756 0.492 0.828 ;
      RECT 0.072 0.252 0.144 0.828 ;
      RECT 1.472 0.252 1.544 0.596 ;
      RECT 0.072 0.252 1.544 0.324 ;
      RECT 0.16 0.108 1.136 0.18 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END MAJ_x2_75t

MACRO MAJ_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MAJ_x3_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.424 0.36 0.656 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.756 1.332 0.828 ;
        RECT 1.26 0.424 1.332 0.828 ;
        RECT 1.132 0.504 1.332 0.576 ;
        RECT 0.592 0.504 0.664 0.828 ;
        RECT 0.484 0.504 0.664 0.576 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.764 0.612 1.008 0.684 ;
        RECT 0.936 0.396 1.008 0.684 ;
        RECT 0.764 0.396 1.008 0.468 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.9 2.016 0.972 ;
        RECT 1.456 0.108 2.016 0.18 ;
        RECT 1.8 0.108 1.872 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.756 0.492 0.828 ;
      RECT 0.072 0.252 0.144 0.828 ;
      RECT 1.472 0.252 1.544 0.596 ;
      RECT 0.072 0.252 1.544 0.324 ;
      RECT 0.16 0.108 1.136 0.18 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END MAJ_x3_75t

MACRO MUX2_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2_x1_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.316 2.304 0.756 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.944 0.304 2.016 0.74 ;
    END
  END B
  PIN O
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.144 0.36 0.216 0.812 ;
        RECT 0.072 0.108 0.144 0.432 ;
    END
  END O
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.484 0.432 1.524 0.504 ;
      LAYER M1 ;
        RECT 1.432 0.412 1.504 0.596 ;
        RECT 0.504 0.268 0.576 0.668 ;
      LAYER V1 ;
        RECT 0.504 0.432 0.576 0.504 ;
        RECT 1.432 0.432 1.504 0.504 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 2.32 0.9 2.52 0.972 ;
      RECT 2.448 0.144 2.52 0.972 ;
      RECT 2.32 0.144 2.52 0.216 ;
      RECT 1.8 0.864 2.036 0.936 ;
      RECT 1.8 0.108 1.872 0.936 ;
      RECT 1.456 0.108 2 0.18 ;
      RECT 1.492 0.72 1.64 0.792 ;
      RECT 1.26 0.34 1.332 0.812 ;
      RECT 1.024 0.144 1.172 0.216 ;
      RECT 1.088 0.484 1.16 0.668 ;
      RECT 0.988 0.864 1.136 0.936 ;
      RECT 0.648 0.184 0.72 0.9 ;
      RECT 0.288 0.484 0.36 0.812 ;
    LAYER M2 ;
      RECT 1.492 0.72 2.54 0.792 ;
      RECT 1.024 0.144 2.432 0.216 ;
      RECT 1.024 0.864 2 0.936 ;
      RECT 0.268 0.72 1.352 0.792 ;
      RECT 0.628 0.576 1.18 0.648 ;
    LAYER V1 ;
      RECT 2.448 0.72 2.52 0.792 ;
      RECT 2.34 0.144 2.412 0.216 ;
      RECT 1.908 0.864 1.98 0.936 ;
      RECT 1.512 0.72 1.584 0.792 ;
      RECT 1.26 0.72 1.332 0.792 ;
      RECT 1.088 0.576 1.16 0.648 ;
      RECT 1.044 0.144 1.116 0.216 ;
      RECT 1.044 0.864 1.116 0.936 ;
      RECT 0.648 0.576 0.72 0.648 ;
      RECT 0.288 0.72 0.36 0.792 ;
  END
END MUX2_x1_75t

MACRO MUX2_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2_x2_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.504 1.388 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.26 1.872 0.596 ;
        RECT 1.724 0.26 1.872 0.332 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Z
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.9 0.704 0.972 ;
        RECT 0.504 0.108 0.704 0.18 ;
        RECT 0.504 0.108 0.576 0.972 ;
    END
  END Z
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.268 0.432 2.172 0.504 ;
      LAYER M1 ;
        RECT 2.08 0.376 2.152 0.596 ;
        RECT 0.288 0.304 0.36 0.776 ;
      LAYER V1 ;
        RECT 0.288 0.432 0.36 0.504 ;
        RECT 2.08 0.432 2.152 0.504 ;
    END
  END S
  OBS
    LAYER M1 ;
      RECT 1.888 0.72 2.304 0.792 ;
      RECT 2.232 0.108 2.304 0.792 ;
      RECT 1.24 0.108 2.304 0.18 ;
      RECT 1.472 0.72 1.656 0.792 ;
      RECT 1.584 0.484 1.656 0.792 ;
      RECT 0.072 0.9 0.272 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.072 0.108 0.272 0.18 ;
      RECT 1.24 0.9 2.216 0.972 ;
      RECT 0.72 0.304 0.792 0.776 ;
    LAYER M2 ;
      RECT 0.7 0.576 2.324 0.648 ;
      RECT 0.052 0.72 1.584 0.792 ;
    LAYER V1 ;
      RECT 2.232 0.576 2.304 0.648 ;
      RECT 1.492 0.72 1.564 0.792 ;
      RECT 0.72 0.576 0.792 0.648 ;
      RECT 0.072 0.72 0.144 0.792 ;
  END
END MUX2_x2_75t

MACRO NAND2_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_x1_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.232 0.972 ;
        RECT 0.072 0.28 0.232 0.352 ;
        RECT 0.072 0.28 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.728 1.008 0.8 ;
        RECT 0.936 0.404 1.008 0.8 ;
        RECT 0.808 0.404 1.008 0.476 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.224 0.972 ;
        RECT 1.152 0.252 1.224 0.972 ;
        RECT 0.808 0.252 1.224 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END NAND2_x1_75t

MACRO NAND2_x1p5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_x1p5_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.896 0.22 0.968 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.968 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 1.028 0.576 ;
        RECT 0.504 0.748 0.652 0.82 ;
        RECT 0.504 0.26 0.652 0.332 ;
        RECT 0.504 0.26 0.576 0.82 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 1.044 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.252 1.352 0.324 ;
      RECT 0.376 0.108 0.9 0.18 ;
  END
END NAND2_x1p5_75t

MACRO NAND2_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_x2_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.94 0.756 1.088 0.828 ;
        RECT 1.016 0.424 1.088 0.828 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.396 1.872 0.708 ;
        RECT 1.288 0.396 1.872 0.468 ;
        RECT 1.288 0.252 1.36 0.468 ;
        RECT 0.8 0.252 1.36 0.324 ;
        RECT 0.288 0.396 0.872 0.468 ;
        RECT 0.8 0.252 0.872 0.468 ;
        RECT 0.288 0.756 0.436 0.828 ;
        RECT 0.288 0.396 0.36 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 2.088 0.972 ;
        RECT 2.016 0.252 2.088 0.972 ;
        RECT 1.672 0.252 2.088 0.324 ;
        RECT 0.072 0.252 0.488 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 2 0.18 ;
  END
END NAND2_x2_75t

MACRO NAND2_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_xp33_75t 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.572 0.108 0.792 0.18 ;
    END
  END Y
END NAND2_xp33_75t

MACRO NAND2_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_xp5_75t 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.424 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.572 0.108 0.792 0.18 ;
    END
  END Y
END NAND2_xp5_75t

MACRO NAND2_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_xp67_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.5 0.38 0.572 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.252 0.22 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 0.812 0.576 ;
        RECT 0.504 0.728 0.648 0.8 ;
        RECT 0.504 0.28 0.648 0.352 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.9 1.224 0.972 ;
        RECT 1.152 0.252 1.224 0.972 ;
        RECT 0.808 0.252 1.224 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END NAND2_xp67_75t

MACRO NAND3_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_x1_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.596 0.756 1.872 0.828 ;
        RECT 1.8 0.424 1.872 0.828 ;
        RECT 1.6 0.424 1.872 0.496 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.972 0.756 1.224 0.828 ;
        RECT 1.152 0.396 1.224 0.828 ;
        RECT 0.984 0.396 1.224 0.468 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.892 0.22 0.964 ;
        RECT 0.072 0.28 0.22 0.352 ;
        RECT 0.072 0.28 0.144 0.964 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 2.304 0.972 ;
        RECT 2.232 0.252 2.304 0.972 ;
        RECT 1.672 0.252 2.304 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.024 0.108 2 0.18 ;
      RECT 0.376 0.252 1.352 0.324 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END NAND3_x1_75t

MACRO NAND3_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_x2_75t 0 0 ;
  SIZE 4.32 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.352 0.756 2.972 0.828 ;
        RECT 2.9 0.424 2.972 0.828 ;
        RECT 1.352 0.424 1.424 0.828 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.188 0.424 2.26 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.32 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 4.248 0.972 ;
        RECT 4.176 0.252 4.248 0.972 ;
        RECT 3.616 0.252 4.248 0.324 ;
        RECT 0.072 0.252 0.704 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.676 0.72 3.632 0.792 ;
      LAYER M1 ;
        RECT 3.464 0.756 3.612 0.828 ;
        RECT 3.54 0.432 3.612 0.828 ;
        RECT 0.696 0.756 0.844 0.828 ;
        RECT 0.696 0.424 0.768 0.828 ;
      LAYER V1 ;
        RECT 0.696 0.72 0.768 0.792 ;
        RECT 3.54 0.72 3.612 0.792 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 2.968 0.108 3.944 0.18 ;
      RECT 1.024 0.252 3.296 0.324 ;
      RECT 1.672 0.108 2.648 0.18 ;
      RECT 0.376 0.108 1.352 0.18 ;
  END
END NAND3_x2_75t

MACRO NAND3_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_xp33_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.728 0.364 0.8 ;
        RECT 0.216 0.28 0.364 0.352 ;
        RECT 0.216 0.28 0.288 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.112 0.576 0.8 ;
        RECT 0.428 0.112 0.576 0.184 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.716 0.728 0.864 0.8 ;
        RECT 0.792 0.136 0.864 0.8 ;
        RECT 0.716 0.136 0.864 0.208 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.704 0.972 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
END NAND3_xp33_75t

MACRO NAND4_xp25_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_xp25_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.108 0.792 0.8 ;
        RECT 0.644 0.108 0.792 0.18 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.728 0.576 0.8 ;
        RECT 0.504 0.284 0.576 0.8 ;
        RECT 0.428 0.284 0.576 0.356 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.728 0.22 0.8 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.8 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.16 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 1.024 0.108 1.224 0.18 ;
    END
  END Y
END NAND4_xp25_75t

MACRO NAND4_xp75_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_xp75_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.588 0.728 2.736 0.8 ;
        RECT 2.664 0.424 2.736 0.8 ;
        RECT 2.588 0.424 2.736 0.496 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.404 2.196 0.476 ;
        RECT 2.124 0.28 2.196 0.476 ;
        RECT 1.8 0.728 1.948 0.8 ;
        RECT 1.8 0.404 1.872 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.86 0.728 1.008 0.8 ;
        RECT 0.936 0.404 1.008 0.8 ;
        RECT 0.828 0.404 1.008 0.476 ;
        RECT 0.828 0.28 0.9 0.476 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.228 0.972 ;
        RECT 0.072 0.108 0.228 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 2.952 0.972 ;
        RECT 2.88 0.252 2.952 0.972 ;
        RECT 2.32 0.252 2.952 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.648 0.108 2.664 0.18 ;
      RECT 1.024 0.252 1.996 0.324 ;
      RECT 0.368 0.108 1.36 0.18 ;
  END
END NAND4_xp75_75t

MACRO NAND5_xp2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND5_xp2_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.212 0.62 0.36 0.692 ;
        RECT 0.288 0.28 0.36 0.692 ;
        RECT 0.212 0.28 0.36 0.352 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.136 0.576 0.828 ;
        RECT 0.428 0.136 0.576 0.208 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.136 0.912 0.208 ;
        RECT 0.72 0.136 0.792 0.8 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.036 0.324 1.228 0.396 ;
        RECT 0.944 0.728 1.108 0.8 ;
        RECT 1.036 0.324 1.108 0.8 ;
        RECT 0.944 0.5 1.108 0.572 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.296 0.728 1.444 0.8 ;
        RECT 1.372 0.136 1.444 0.8 ;
        RECT 1.22 0.5 1.444 0.572 ;
        RECT 1.296 0.136 1.444 0.208 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.036 0.9 1.444 0.972 ;
        RECT 0.036 0.108 0.28 0.18 ;
        RECT 0.036 0.108 0.108 0.972 ;
    END
  END Y
END NAND5_xp2_75t

MACRO NOR2_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_x1_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 0.92 0.576 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.376 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END NOR2_x1_75t

MACRO NOR2_x1p5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_x1p5_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.336 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 1.028 0.576 ;
        RECT 0.504 0.252 0.652 0.324 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.376 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.756 1.352 0.828 ;
      RECT 0.376 0.9 0.9 0.972 ;
  END
END NOR2_x1p5_75t

MACRO NOR2_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_x2_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.656 ;
        RECT 0.86 0.252 1.008 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.288 0.612 1.872 0.684 ;
        RECT 1.8 0.372 1.872 0.684 ;
        RECT 0.72 0.756 1.36 0.828 ;
        RECT 1.288 0.612 1.36 0.828 ;
        RECT 0.72 0.612 0.792 0.828 ;
        RECT 0.288 0.612 0.792 0.684 ;
        RECT 0.288 0.252 0.436 0.324 ;
        RECT 0.288 0.252 0.36 0.684 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.756 2.088 0.828 ;
        RECT 2.016 0.108 2.088 0.828 ;
        RECT 0.072 0.108 2.088 0.18 ;
        RECT 0.072 0.756 0.488 0.828 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 2 0.972 ;
  END
END NOR2_x2_75t

MACRO NOR2_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_xp33_75t 0 0 ;
  SIZE 0.864 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.864 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.864 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.572 0.9 0.792 0.972 ;
        RECT 0.72 0.108 0.792 0.972 ;
        RECT 0.376 0.108 0.792 0.18 ;
    END
  END Y
END NOR2_xp33_75t

MACRO NOR2_xp67_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_xp67_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.508 0.38 0.58 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.504 1.028 0.576 ;
        RECT 0.504 0.252 0.652 0.324 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.756 1.224 0.828 ;
        RECT 1.152 0.108 1.224 0.828 ;
        RECT 0.592 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END NOR2_xp67_75t

MACRO NOR3_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_x1_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.612 1.872 0.684 ;
        RECT 1.8 0.252 1.872 0.684 ;
        RECT 1.584 0.252 1.872 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.612 1.224 0.684 ;
        RECT 1.152 0.252 1.224 0.684 ;
        RECT 0.936 0.252 1.224 0.324 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.36 0.576 ;
        RECT 0.072 0.756 0.22 0.828 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.672 0.756 2.304 0.828 ;
        RECT 2.232 0.108 2.304 0.828 ;
        RECT 0.808 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.024 0.9 2 0.972 ;
      RECT 0.376 0.756 1.352 0.828 ;
      RECT 0.16 0.9 0.704 0.972 ;
  END
END NOR3_x1_75t

MACRO NOR3_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_x2_75t 0 0 ;
  SIZE 4.32 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.9 0.252 2.972 0.656 ;
        RECT 1.368 0.252 2.972 0.324 ;
        RECT 1.368 0.252 1.44 0.656 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.94 0.612 2.596 0.684 ;
        RECT 1.94 0.396 2.596 0.468 ;
        RECT 2.232 0.396 2.304 0.684 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 4.32 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 4.32 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 3.616 0.756 4.248 0.828 ;
        RECT 4.176 0.108 4.248 0.828 ;
        RECT 0.072 0.108 4.248 0.18 ;
        RECT 0.072 0.756 0.704 0.828 ;
        RECT 0.072 0.108 0.144 0.828 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.484 0.288 3.62 0.36 ;
      LAYER M1 ;
        RECT 3.528 0.252 3.6 0.648 ;
        RECT 3.452 0.252 3.6 0.324 ;
        RECT 0.504 0.252 0.652 0.324 ;
        RECT 0.504 0.252 0.576 0.656 ;
      LAYER V1 ;
        RECT 0.504 0.288 0.576 0.36 ;
        RECT 3.528 0.288 3.6 0.36 ;
    END
  END A
  OBS
    LAYER M1 ;
      RECT 2.968 0.9 3.944 0.972 ;
      RECT 1.024 0.756 3.296 0.828 ;
      RECT 1.672 0.9 2.648 0.972 ;
      RECT 0.376 0.9 1.352 0.972 ;
  END
END NOR3_x2_75t

MACRO NOR3_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_xp33_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.224 0.728 0.372 0.8 ;
        RECT 0.224 0.252 0.372 0.324 ;
        RECT 0.224 0.252 0.296 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.9 0.652 0.972 ;
        RECT 0.504 0.396 0.652 0.468 ;
        RECT 0.504 0.396 0.576 0.972 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.792 0.872 0.94 0.944 ;
        RECT 0.792 0.28 0.94 0.352 ;
        RECT 0.792 0.28 0.864 0.944 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.004 0.108 0.684 0.18 ;
        RECT 0.004 0.9 0.252 0.972 ;
        RECT 0.004 0.108 0.076 0.972 ;
    END
  END Y
END NOR3_xp33_75t

MACRO NOR4_xp25_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_xp25_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.252 1.008 0.8 ;
        RECT 0.716 0.252 1.008 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.872 0.868 0.944 ;
        RECT 0.72 0.44 0.792 0.944 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.872 0.576 0.944 ;
        RECT 0.504 0.28 0.576 0.944 ;
        RECT 0.428 0.28 0.576 0.352 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.14 0.872 0.288 0.944 ;
        RECT 0.216 0.28 0.288 0.944 ;
        RECT 0.14 0.28 0.288 0.352 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.16 0.108 1.224 0.18 ;
    END
  END Y
END NOR4_xp25_75t

MACRO NOR4_xp75_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_xp75_75t 0 0 ;
  SIZE 3.024 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.444 0.612 2.736 0.684 ;
        RECT 2.664 0.252 2.736 0.684 ;
        RECT 2.444 0.252 2.736 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.124 0.604 2.196 0.8 ;
        RECT 2.016 0.604 2.196 0.676 ;
        RECT 2.016 0.252 2.088 0.676 ;
        RECT 1.94 0.252 2.088 0.324 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.604 1.224 0.676 ;
        RECT 1.152 0.252 1.224 0.676 ;
        RECT 1.076 0.252 1.224 0.324 ;
        RECT 0.828 0.604 0.9 0.8 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.228 0.972 ;
        RECT 0.072 0.108 0.228 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.024 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.024 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.32 0.756 2.952 0.828 ;
        RECT 2.88 0.108 2.952 0.828 ;
        RECT 0.376 0.108 2.952 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.648 0.9 2.664 0.972 ;
      RECT 1.024 0.756 1.996 0.828 ;
      RECT 0.368 0.9 1.36 0.972 ;
  END
END NOR4_xp75_75t

MACRO NOR5_xp2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR5_xp2_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.212 0.872 0.36 0.944 ;
        RECT 0.288 0.416 0.36 0.944 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.252 0.576 0.944 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.9 1.084 0.972 ;
        RECT 0.72 0.252 0.868 0.324 ;
        RECT 0.72 0.252 0.792 0.972 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.728 1.084 0.8 ;
        RECT 0.936 0.384 1.008 0.8 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.328 1.44 0.944 ;
        RECT 1.148 0.508 1.44 0.58 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 1.352 0.18 ;
        RECT 0.072 0.108 0.144 0.744 ;
    END
  END Y
END NOR5_xp2_75t

MACRO O2A1O1I_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN O2A1O1I_xp33_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.728 0.576 0.8 ;
        RECT 0.504 0.424 0.576 0.8 ;
        RECT 0.428 0.424 0.576 0.496 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1 0.728 0.292 0.8 ;
        RECT 0.22 0.424 0.292 0.8 ;
        RECT 0.1 0.424 0.292 0.496 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.728 0.812 0.8 ;
        RECT 0.648 0.504 0.812 0.576 ;
        RECT 0.648 0.504 0.72 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.824 ;
        RECT 0.828 0.28 1.008 0.352 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 0.376 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.9 0.972 ;
      RECT 0.16 0.252 0.704 0.324 ;
  END
END O2A1O1I_xp33_75t

MACRO O2A1O1I_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN O2A1O1I_xp5_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.052 0.432 1.028 0.504 ;
      LAYER M1 ;
        RECT 0.936 0.412 1.008 0.596 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
      LAYER V1 ;
        RECT 0.072 0.432 0.144 0.504 ;
        RECT 0.936 0.432 1.008 0.504 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.26 0.576 0.656 ;
        RECT 0.364 0.26 0.576 0.332 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.252 1.224 0.656 ;
        RECT 1.076 0.252 1.224 0.324 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.44 0.252 1.512 0.656 ;
        RECT 1.364 0.252 1.512 0.324 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 1.26 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.504 0.756 1.352 0.828 ;
      RECT 0.592 0.108 1.116 0.18 ;
      RECT 0.376 0.9 0.92 0.972 ;
  END
END O2A1O1I_xp5_75t

MACRO OA211_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211_x1_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.344 0.756 0.576 0.828 ;
        RECT 0.504 0.396 0.576 0.828 ;
        RECT 0.428 0.396 0.576 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.748 0.22 0.82 ;
        RECT 0.072 0.26 0.22 0.332 ;
        RECT 0.072 0.26 0.144 0.82 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.748 0.868 0.82 ;
        RECT 0.72 0.424 0.792 0.82 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.404 1.084 0.476 ;
        RECT 0.936 0.404 1.008 0.656 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.22 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.144 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.116 0.972 ;
      RECT 1.044 0.736 1.116 0.972 ;
      RECT 1.044 0.736 1.28 0.808 ;
      RECT 1.208 0.252 1.28 0.808 ;
      RECT 0.396 0.252 1.28 0.324 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END OA211_x1_75t

MACRO OA211_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA211_x2_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.348 0.748 0.576 0.82 ;
        RECT 0.504 0.404 0.576 0.82 ;
        RECT 0.424 0.404 0.576 0.476 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.748 0.224 0.82 ;
        RECT 0.072 0.26 0.224 0.332 ;
        RECT 0.072 0.26 0.144 0.82 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.748 0.872 0.82 ;
        RECT 0.72 0.424 0.792 0.82 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.604 1.16 0.676 ;
        RECT 0.936 0.404 1.16 0.476 ;
        RECT 0.936 0.404 1.008 0.676 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.24 0.9 1.584 0.972 ;
        RECT 1.512 0.108 1.584 0.972 ;
        RECT 1.144 0.108 1.584 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 1.116 0.972 ;
      RECT 1.044 0.756 1.116 0.972 ;
      RECT 1.044 0.756 1.44 0.828 ;
      RECT 1.368 0.252 1.44 0.828 ;
      RECT 0.396 0.252 1.44 0.324 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END OA211_x2_75t

MACRO OA21_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21_x2_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.26 0.22 0.332 ;
        RECT 0.072 0.26 0.144 0.972 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.504 0.596 0.576 ;
        RECT 0.288 0.752 0.436 0.824 ;
        RECT 0.288 0.424 0.36 0.824 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.612 0.956 0.684 ;
        RECT 0.72 0.424 0.792 0.684 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.024 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.592 0.9 0.896 0.972 ;
      RECT 0.824 0.756 0.896 0.972 ;
      RECT 0.824 0.756 1.224 0.828 ;
      RECT 1.152 0.252 1.224 0.828 ;
      RECT 0.396 0.252 1.224 0.324 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END OA21_x2_75t

MACRO OA221_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221_x1_75t 0 0 ;
  SIZE 3.24 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.756 0.836 0.828 ;
        RECT 0.504 0.396 0.836 0.468 ;
        RECT 0.504 0.396 0.576 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.756 1.376 0.828 ;
        RECT 0.936 0.396 1.376 0.468 ;
        RECT 0.936 0.396 1.008 0.828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.972 0.756 2.304 0.828 ;
        RECT 2.232 0.396 2.304 0.828 ;
        RECT 1.972 0.396 2.304 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.5 0.756 1.872 0.828 ;
        RECT 1.8 0.396 1.872 0.828 ;
        RECT 1.5 0.396 1.872 0.468 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.664 0.756 2.996 0.828 ;
        RECT 2.664 0.396 2.996 0.468 ;
        RECT 2.664 0.396 2.736 0.828 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.24 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.068 0.108 0.272 0.18 ;
        RECT 0.124 0.576 0.196 0.832 ;
        RECT 0.068 0.108 0.14 0.648 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.288 0.9 3.168 0.972 ;
      RECT 3.096 0.252 3.168 0.972 ;
      RECT 0.288 0.484 0.36 0.972 ;
      RECT 2.748 0.252 3.168 0.324 ;
      RECT 1.672 0.108 3.08 0.18 ;
      RECT 0.592 0.252 2.456 0.324 ;
  END
END OA221_x1_75t

MACRO OA221_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA221_x2_75t 0 0 ;
  SIZE 3.456 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.748 0.756 1.008 0.828 ;
        RECT 0.936 0.396 1.008 0.828 ;
        RECT 0.748 0.396 1.008 0.468 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.108 0.756 1.628 0.828 ;
        RECT 1.108 0.396 1.628 0.468 ;
        RECT 1.368 0.396 1.44 0.828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.188 0.756 2.52 0.828 ;
        RECT 2.448 0.396 2.52 0.828 ;
        RECT 2.188 0.396 2.52 0.468 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.752 0.756 2.088 0.828 ;
        RECT 2.016 0.396 2.088 0.828 ;
        RECT 1.752 0.396 2.088 0.468 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.62 0.756 3.212 0.828 ;
        RECT 2.62 0.396 3.212 0.468 ;
        RECT 2.88 0.396 2.952 0.828 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.456 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.456 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.9 0.468 0.972 ;
        RECT 0.396 0.756 0.468 0.972 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.576 0.9 3.384 0.972 ;
      RECT 3.312 0.252 3.384 0.972 ;
      RECT 0.576 0.504 0.648 0.972 ;
      RECT 0.484 0.504 0.648 0.576 ;
      RECT 2.964 0.252 3.384 0.324 ;
      RECT 1.888 0.108 3.296 0.18 ;
      RECT 0.808 0.252 2.672 0.324 ;
  END
END OA221_x2_75t

MACRO OA222_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222_x1_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.244 0.756 0.404 0.828 ;
        RECT 0.244 0.396 0.404 0.468 ;
        RECT 0.288 0.396 0.36 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.004 0.756 1.152 0.828 ;
        RECT 1.004 0.396 1.152 0.468 ;
        RECT 1.004 0.396 1.076 0.828 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.756 0.904 0.828 ;
        RECT 0.72 0.396 0.904 0.468 ;
        RECT 0.72 0.396 0.792 0.828 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.276 0.756 1.656 0.828 ;
        RECT 1.584 0.28 1.656 0.828 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 2.108 0.352 ;
        RECT 1.756 0.756 1.916 0.828 ;
        RECT 1.8 0.28 1.872 0.828 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.108 2.304 0.54 ;
        RECT 2.16 0.468 2.232 0.8 ;
        RECT 2.104 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 2.088 0.972 ;
      RECT 2.016 0.484 2.088 0.972 ;
      RECT 0.072 0.252 0.144 0.972 ;
      RECT 0.072 0.252 0.488 0.324 ;
      RECT 0.808 0.252 1.44 0.324 ;
      RECT 1.368 0.108 1.44 0.324 ;
      RECT 1.368 0.108 1.872 0.18 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END OA222_x1_75t

MACRO OA222_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA222_x2_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.756 0.404 0.828 ;
        RECT 0.216 0.396 0.404 0.468 ;
        RECT 0.216 0.396 0.288 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.004 0.756 1.304 0.828 ;
        RECT 1.004 0.396 1.304 0.468 ;
        RECT 1.004 0.396 1.076 0.828 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.756 0.904 0.828 ;
        RECT 0.72 0.396 0.904 0.468 ;
        RECT 0.72 0.396 0.792 0.828 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.428 0.756 1.656 0.828 ;
        RECT 1.584 0.28 1.656 0.828 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 2.348 0.352 ;
        RECT 1.8 0.28 1.872 0.8 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.124 0.9 2.52 0.972 ;
        RECT 2.448 0.108 2.52 0.972 ;
        RECT 2.104 0.108 2.52 0.18 ;
        RECT 2.124 0.676 2.196 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 2.016 0.972 ;
      RECT 1.944 0.504 2.016 0.972 ;
      RECT 0.072 0.252 0.144 0.972 ;
      RECT 1.944 0.504 2.216 0.576 ;
      RECT 0.072 0.252 0.488 0.324 ;
      RECT 0.808 0.252 1.44 0.324 ;
      RECT 1.368 0.108 1.44 0.324 ;
      RECT 1.368 0.108 1.872 0.18 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END OA222_x2_75t

MACRO OA22_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22_x2_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.756 1.152 0.828 ;
        RECT 1.08 0.424 1.152 0.828 ;
        RECT 0.936 0.424 1.008 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.252 0.756 1.44 0.828 ;
        RECT 1.368 0.424 1.44 0.828 ;
        RECT 1.252 0.424 1.44 0.496 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.9 2.012 0.972 ;
        RECT 1.8 0.252 2.012 0.324 ;
        RECT 1.8 0.252 1.872 0.972 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.252 1.656 0.8 ;
        RECT 1.508 0.252 1.656 0.324 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.488 0.972 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.72 0.9 1.568 0.972 ;
      RECT 0.72 0.252 0.792 0.972 ;
      RECT 0.504 0.504 0.792 0.576 ;
      RECT 0.72 0.252 1.332 0.324 ;
      RECT 1.024 0.108 2 0.18 ;
  END
END OA22_x2_75t

MACRO OA31_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA31_x2_75t 0 0 ;
  SIZE 3.24 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.756 0.404 0.828 ;
        RECT 0.216 0.396 0.404 0.468 ;
        RECT 0.216 0.396 0.288 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.396 1.008 0.656 ;
        RECT 0.504 0.396 1.008 0.468 ;
        RECT 0.504 0.756 0.684 0.828 ;
        RECT 0.504 0.396 0.576 0.828 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.504 1.656 0.576 ;
        RECT 1.368 0.252 1.44 0.656 ;
        RECT 1.292 0.252 1.44 0.324 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.404 2.308 0.476 ;
        RECT 1.796 0.612 2.088 0.684 ;
        RECT 2.016 0.404 2.088 0.684 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 3.24 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 3.24 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.772 0.9 3.168 0.972 ;
        RECT 3.096 0.108 3.168 0.972 ;
        RECT 2.772 0.108 3.168 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.476 0.756 2.52 0.828 ;
      RECT 2.448 0.252 2.52 0.828 ;
      RECT 2.448 0.504 2.668 0.576 ;
      RECT 1.672 0.252 2.52 0.324 ;
      RECT 1.268 0.9 1.784 0.972 ;
      RECT 1.268 0.756 1.34 0.972 ;
      RECT 0.808 0.756 1.34 0.828 ;
      RECT 0.376 0.108 2 0.18 ;
      RECT 0.16 0.252 1.136 0.324 ;
      RECT 0.16 0.9 1.136 0.972 ;
  END
END OA31_x2_75t

MACRO OA331_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA331_x1_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.62 0.728 0.792 0.8 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.624 ;
        RECT 0.404 0.28 0.576 0.352 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.144 0.424 1.216 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.756 1.756 0.828 ;
        RECT 1.584 0.424 1.656 0.828 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.672 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.9 2.088 0.972 ;
      RECT 2.016 0.108 2.088 0.972 ;
      RECT 0.396 0.744 0.468 0.972 ;
      RECT 0.288 0.744 0.468 0.816 ;
      RECT 0.288 0.46 0.36 0.816 ;
      RECT 1.908 0.108 2.088 0.18 ;
      RECT 0.936 0.252 1.572 0.324 ;
      RECT 0.936 0.108 1.008 0.324 ;
      RECT 0.592 0.108 1.008 0.18 ;
      RECT 1.232 0.108 1.764 0.18 ;
  END
END OA331_x1_75t

MACRO OA331_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA331_x2_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.076 0.756 1.224 0.828 ;
        RECT 1.152 0.424 1.224 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.664 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.664 ;
        RECT 0.384 0.28 0.792 0.352 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.756 1.732 0.828 ;
        RECT 1.584 0.424 1.656 0.828 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.424 1.872 0.708 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.424 2.164 0.496 ;
        RECT 2.016 0.424 2.088 0.768 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.9 0.488 0.972 ;
        RECT 0.18 0.108 0.488 0.18 ;
        RECT 0.18 0.108 0.252 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.9 2.304 0.972 ;
      RECT 2.232 0.796 2.304 0.972 ;
      RECT 0.612 0.744 0.684 0.972 ;
      RECT 0.504 0.744 0.684 0.816 ;
      RECT 0.504 0.46 0.576 0.816 ;
      RECT 1.152 0.252 1.788 0.324 ;
      RECT 1.152 0.108 1.224 0.324 ;
      RECT 0.808 0.108 1.224 0.18 ;
      RECT 2.156 0.252 2.304 0.324 ;
      RECT 1.448 0.108 2.004 0.18 ;
  END
END OA331_x2_75t

MACRO OA332_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA332_x1_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.424 1.656 0.8 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.076 0.424 2.148 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.824 0.424 1.896 0.8 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.376 0.972 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.504 0.9 2.304 0.972 ;
      RECT 2.232 0.252 2.304 0.972 ;
      RECT 0.504 0.756 0.576 0.972 ;
      RECT 0.288 0.756 0.576 0.828 ;
      RECT 0.288 0.28 0.36 0.828 ;
      RECT 1.884 0.252 2.304 0.324 ;
      RECT 0.936 0.252 1.548 0.324 ;
      RECT 0.936 0.108 1.008 0.324 ;
      RECT 0.584 0.108 1.008 0.18 ;
      RECT 1.232 0.108 2.224 0.18 ;
  END
END OA332_x1_75t

MACRO OA332_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA332_x2_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.424 1.656 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.424 1.872 0.8 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.424 2.304 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.424 2.088 0.8 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.548 0.972 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.72 0.9 2.52 0.972 ;
      RECT 2.448 0.252 2.52 0.972 ;
      RECT 0.72 0.756 0.792 0.972 ;
      RECT 0.504 0.756 0.792 0.828 ;
      RECT 0.504 0.476 0.576 0.828 ;
      RECT 2.1 0.252 2.52 0.324 ;
      RECT 1.152 0.252 1.788 0.324 ;
      RECT 1.152 0.108 1.224 0.324 ;
      RECT 0.8 0.108 1.224 0.18 ;
      RECT 1.448 0.108 2.44 0.18 ;
  END
END OA332_x2_75t

MACRO OA333_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA333_x1_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.424 2.304 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.424 2.088 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.424 1.872 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.424 1.656 0.8 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.656 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.9 2.52 0.972 ;
      RECT 2.448 0.252 2.52 0.972 ;
      RECT 0.396 0.744 0.468 0.972 ;
      RECT 0.288 0.744 0.468 0.816 ;
      RECT 0.288 0.46 0.36 0.816 ;
      RECT 1.868 0.252 2.52 0.324 ;
      RECT 0.928 0.252 1.576 0.324 ;
      RECT 0.928 0.108 1 0.324 ;
      RECT 0.588 0.108 1 0.18 ;
      RECT 1.236 0.108 2.276 0.18 ;
  END
END OA333_x1_75t

MACRO OA333_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA333_x2_75t 0 0 ;
  SIZE 2.808 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.448 0.424 2.52 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.232 0.424 2.304 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0.424 2.088 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.424 1.656 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.424 1.872 0.8 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.656 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.808 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.808 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.9 0.488 0.972 ;
        RECT 0.288 0.108 0.488 0.18 ;
        RECT 0.288 0.108 0.36 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.9 2.736 0.972 ;
      RECT 2.664 0.252 2.736 0.972 ;
      RECT 0.612 0.744 0.684 0.972 ;
      RECT 0.504 0.744 0.684 0.816 ;
      RECT 0.504 0.46 0.576 0.816 ;
      RECT 2.084 0.252 2.736 0.324 ;
      RECT 1.144 0.252 1.792 0.324 ;
      RECT 1.144 0.108 1.216 0.324 ;
      RECT 0.804 0.108 1.216 0.18 ;
      RECT 1.452 0.108 2.492 0.18 ;
  END
END OA333_x2_75t

MACRO OA33_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA33_x2_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.316 0.792 0.656 ;
        RECT 0.288 0.316 0.792 0.388 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.748 0.756 1.008 0.828 ;
        RECT 0.936 0.404 1.008 0.828 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.252 1.224 0.8 ;
        RECT 1.076 0.252 1.224 0.324 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.756 1.948 0.828 ;
        RECT 1.8 0.396 1.948 0.468 ;
        RECT 1.8 0.396 1.872 0.828 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.424 1.656 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.9 0.468 0.972 ;
        RECT 0.396 0.808 0.468 0.972 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.576 0.9 2.12 0.972 ;
      RECT 2.048 0.252 2.12 0.972 ;
      RECT 0.576 0.504 0.648 0.972 ;
      RECT 0.484 0.504 0.648 0.576 ;
      RECT 1.456 0.252 2.12 0.324 ;
      RECT 0.808 0.108 1.784 0.18 ;
  END
END OA33_x2_75t

MACRO OAI211_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211_x1_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.784 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.204 0.576 1.028 0.648 ;
      LAYER M1 ;
        RECT 0.936 0.48 1.008 0.664 ;
        RECT 0.224 0.428 0.296 0.684 ;
      LAYER V1 ;
        RECT 0.224 0.576 0.296 0.648 ;
        RECT 0.936 0.576 1.008 0.648 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.132 0.432 1.892 0.504 ;
      LAYER M1 ;
        RECT 1.8 0.412 1.872 0.664 ;
        RECT 1.152 0.412 1.224 0.78 ;
      LAYER V1 ;
        RECT 1.152 0.432 1.224 0.504 ;
        RECT 1.8 0.432 1.872 0.504 ;
    END
  END B
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.164 0.864 2 0.936 ;
      LAYER M1 ;
        RECT 1.888 0.864 2 0.936 ;
        RECT 1.456 0.864 1.568 0.936 ;
        RECT 1.024 0.864 1.136 0.936 ;
        RECT 0.072 0.252 0.884 0.324 ;
        RECT 0.072 0.864 0.256 0.936 ;
        RECT 0.072 0.252 0.144 0.936 ;
      LAYER V1 ;
        RECT 0.164 0.864 0.236 0.936 ;
        RECT 1.044 0.864 1.116 0.936 ;
        RECT 1.476 0.864 1.548 0.936 ;
        RECT 1.908 0.864 1.98 0.936 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.108 1.116 0.292 ;
      RECT 0.16 0.108 1.116 0.18 ;
      RECT 0.396 0.9 0.9 0.972 ;
      RECT 0.828 0.788 0.9 0.972 ;
      RECT 1.908 0.144 2.02 0.216 ;
      RECT 1.24 0.108 1.784 0.18 ;
    LAYER M2 ;
      RECT 1.024 0.144 2.02 0.216 ;
    LAYER V1 ;
      RECT 1.928 0.144 2 0.216 ;
      RECT 1.044 0.144 1.116 0.216 ;
  END
END OAI211_x1_75t

MACRO OAI211_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211_xp5_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.748 0.576 0.82 ;
        RECT 0.504 0.424 0.576 0.82 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.36 0.576 ;
        RECT 0.072 0.748 0.22 0.82 ;
        RECT 0.072 0.396 0.144 0.82 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.392 0.792 0.72 ;
        RECT 0.648 0.648 0.72 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.16 0.9 1.152 0.972 ;
        RECT 1.08 0.108 1.152 0.972 ;
        RECT 0.396 0.108 1.152 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.252 0.672 0.324 ;
      RECT 0.18 0.18 0.252 0.324 ;
  END
END OAI211_xp5_75t

MACRO OAI21_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_x1_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.756 1.224 0.828 ;
        RECT 1.152 0.424 1.224 0.828 ;
        RECT 0.504 0.424 0.576 0.828 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.648 0.508 1.024 0.58 ;
        RECT 0.648 0.424 0.72 0.656 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.252 1.44 0.616 ;
        RECT 0.32 0.252 1.44 0.324 ;
        RECT 0.216 0.312 0.392 0.384 ;
        RECT 0.216 0.312 0.288 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 1.476 0.108 1.656 0.18 ;
        RECT 0.072 0.108 0.252 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.108 1.332 0.18 ;
  END
END OAI21_x1_75t

MACRO OAI21_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_xp33_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.86 0.22 0.944 ;
        RECT 0.072 0.252 0.22 0.336 ;
        RECT 0.072 0.252 0.144 0.944 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.284 0.74 0.576 0.812 ;
        RECT 0.504 0.424 0.576 0.812 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.72 ;
        RECT 0.648 0.648 0.72 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.9 1.008 0.972 ;
        RECT 0.936 0.252 1.008 0.972 ;
        RECT 0.396 0.252 1.008 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.108 0.704 0.18 ;
  END
END OAI21_xp33_75t

MACRO OAI21_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_xp5_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.28 0.144 0.944 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.74 0.576 0.812 ;
        RECT 0.504 0.424 0.576 0.812 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.716 0.748 0.864 0.82 ;
        RECT 0.792 0.424 0.864 0.82 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.592 0.9 1.008 0.972 ;
        RECT 0.936 0.252 1.008 0.972 ;
        RECT 0.396 0.252 1.008 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 0.704 0.18 ;
  END
END OAI21_xp5_75t

MACRO OAI221_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221_xp5_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.384 1.008 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.148 0.9 1.44 0.972 ;
        RECT 1.368 0.28 1.44 0.972 ;
        RECT 1.224 0.504 1.44 0.576 ;
        RECT 1.148 0.28 1.44 0.352 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.076 0.728 0.288 0.8 ;
        RECT 0.216 0.28 0.288 0.8 ;
        RECT 0.076 0.28 0.288 0.352 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.384 0.792 0.72 ;
        RECT 0.648 0.648 0.72 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.9 0.92 0.972 ;
        RECT 0.36 0.28 0.432 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.828 0.108 0.9 0.312 ;
      RECT 0.828 0.108 1.352 0.18 ;
      RECT 0.16 0.108 0.684 0.18 ;
  END
END OAI221_xp5_75t

MACRO OAI222_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222_xp33_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.28 0.288 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.728 1.4 0.8 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.74 ;
        RECT 0.648 0.652 0.72 0.8 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.72 ;
        RECT 1.512 0.648 1.584 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.8 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.9 2.088 0.972 ;
        RECT 2.016 0.22 2.088 0.972 ;
        RECT 0.36 0.28 0.432 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.808 0.252 1.44 0.324 ;
      RECT 1.368 0.108 1.44 0.324 ;
      RECT 1.368 0.108 1.872 0.18 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END OAI222_xp33_75t

MACRO OAI22_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_x1_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.612 1.7 0.684 ;
        RECT 1.368 0.396 1.516 0.468 ;
        RECT 1.368 0.396 1.44 0.684 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.756 1.872 0.828 ;
        RECT 1.8 0.396 1.872 0.828 ;
        RECT 1.724 0.396 1.872 0.468 ;
        RECT 1.152 0.404 1.224 0.828 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.572 0.612 0.72 0.684 ;
        RECT 0.648 0.252 0.72 0.684 ;
        RECT 0.572 0.252 0.72 0.324 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.756 1.008 0.828 ;
        RECT 0.936 0.28 1.008 0.828 ;
        RECT 0.216 0.252 0.436 0.324 ;
        RECT 0.216 0.252 0.288 0.828 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.152 0.9 2.088 0.972 ;
        RECT 2.016 0.252 2.088 0.972 ;
        RECT 1.236 0.252 2.088 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 2 0.18 ;
  END
END OAI22_x1_75t

MACRO OAI22_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_xp33_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.424 0.36 0.72 ;
        RECT 0.216 0.648 0.288 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.008 0.9 1.224 0.972 ;
        RECT 1.152 0.28 1.224 0.972 ;
        RECT 1.008 0.504 1.224 0.576 ;
        RECT 1.008 0.28 1.224 0.352 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.72 ;
        RECT 0.648 0.648 0.72 0.8 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.704 0.972 ;
        RECT 0.072 0.252 0.468 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END OAI22_xp33_75t

MACRO OAI22_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_xp5_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.424 0.36 0.72 ;
        RECT 0.216 0.648 0.288 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.404 0.576 0.8 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.008 0.9 1.224 0.972 ;
        RECT 1.152 0.28 1.224 0.972 ;
        RECT 1.008 0.504 1.224 0.576 ;
        RECT 1.008 0.28 1.224 0.352 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.792 0.68 0.864 0.892 ;
        RECT 0.72 0.252 0.792 0.752 ;
        RECT 0.604 0.252 0.792 0.324 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.704 0.972 ;
        RECT 0.072 0.252 0.468 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.108 1.136 0.18 ;
  END
END OAI22_xp5_75t

MACRO OAI311_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI311_xp33_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.812 ;
        RECT 0.648 0.74 0.72 0.892 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.944 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.136 0.144 0.944 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.26 1.008 0.8 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.26 1.224 0.72 ;
        RECT 1.08 0.648 1.152 0.8 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 1.44 0.972 ;
        RECT 1.368 0.108 1.44 0.972 ;
        RECT 1.24 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.108 0.92 0.18 ;
  END
END OAI311_xp33_75t

MACRO OAI31_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31_xp33_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
        RECT 0.648 0.728 0.72 0.88 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.944 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.508 0.288 0.58 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A3
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.804 0.9 1.224 0.972 ;
        RECT 1.152 0.108 1.224 0.972 ;
        RECT 1.044 0.108 1.224 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.372 0.108 0.9 0.18 ;
  END
END OAI31_xp33_75t

MACRO OAI321_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI321_xp33_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.324 0.792 0.808 ;
        RECT 0.648 0.736 0.72 0.888 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.944 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.38 0.576 ;
        RECT 0.072 0.9 0.236 0.972 ;
        RECT 0.072 0.108 0.236 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.404 1.224 0.72 ;
        RECT 1.08 0.648 1.152 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.324 1.008 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.808 0.9 1.656 0.972 ;
        RECT 1.584 0.252 1.656 0.972 ;
        RECT 1.24 0.252 1.656 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.828 0.108 0.9 0.252 ;
      RECT 0.396 0.108 0.9 0.18 ;
      RECT 1.024 0.108 1.584 0.18 ;
  END
END OAI321_xp33_75t

MACRO OAI322_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI322_xp33_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.424 0.792 0.72 ;
        RECT 0.648 0.648 0.72 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.404 1.224 0.72 ;
        RECT 1.08 0.648 1.152 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.748 0.576 0.82 ;
        RECT 0.504 0.404 0.576 0.82 ;
        RECT 0.428 0.404 0.576 0.476 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.288 0.576 ;
        RECT 0.072 0.872 0.228 0.944 ;
        RECT 0.072 0.28 0.228 0.352 ;
        RECT 0.072 0.28 0.144 0.944 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.424 1.656 0.72 ;
        RECT 1.512 0.648 1.584 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.404 1.44 0.8 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.588 0.9 1.872 0.972 ;
        RECT 1.8 0.252 1.872 0.972 ;
        RECT 1.456 0.252 1.872 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.612 0.252 1.136 0.324 ;
      RECT 0.612 0.108 0.684 0.324 ;
      RECT 0.16 0.108 0.684 0.18 ;
      RECT 0.808 0.108 1.8 0.18 ;
  END
END OAI322_xp33_75t

MACRO OAI32_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32_xp33_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.288 0.576 ;
        RECT 0.072 0.728 0.22 0.8 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.252 0.888 0.324 ;
        RECT 0.72 0.252 0.792 0.72 ;
        RECT 0.648 0.648 0.72 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.424 1.008 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.72 ;
        RECT 1.08 0.648 1.152 0.8 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.16 0.9 1.44 0.972 ;
        RECT 1.368 0.252 1.44 0.972 ;
        RECT 1.024 0.252 1.44 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.108 1.352 0.18 ;
  END
END OAI32_xp33_75t

MACRO OAI331_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI331_xp33_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.808 ;
        RECT 0.648 0.736 0.72 0.888 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.9 0.576 0.972 ;
        RECT 0.504 0.28 0.576 0.972 ;
        RECT 0.428 0.28 0.576 0.352 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.288 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.396 1.008 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.72 ;
        RECT 1.08 0.648 1.152 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.656 0.308 1.728 0.476 ;
        RECT 1.584 0.404 1.656 0.72 ;
        RECT 1.512 0.648 1.584 0.8 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.804 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.668 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.252 1.548 0.324 ;
      RECT 1.476 0.16 1.548 0.324 ;
      RECT 0.376 0.108 1.332 0.18 ;
  END
END OAI331_xp33_75t

MACRO OAI332_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI332_xp33_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.796 ;
        RECT 0.648 0.724 0.72 0.876 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.9 0.576 0.972 ;
        RECT 0.504 0.28 0.576 0.972 ;
        RECT 0.428 0.28 0.576 0.352 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.288 0.576 ;
        RECT 0.072 0.9 0.264 0.972 ;
        RECT 0.072 0.108 0.264 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.396 1.008 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.72 ;
        RECT 1.08 0.648 1.152 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.424 1.872 0.8 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.656 0.648 1.728 0.8 ;
        RECT 1.584 0.404 1.656 0.72 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.804 0.9 2.088 0.972 ;
        RECT 2.016 0.252 2.088 0.972 ;
        RECT 1.692 0.252 2.088 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.252 1.548 0.324 ;
      RECT 1.476 0.108 1.548 0.324 ;
      RECT 1.476 0.108 2.008 0.18 ;
      RECT 0.396 0.108 1.332 0.18 ;
  END
END OAI332_xp33_75t

MACRO OAI333_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI333_xp33_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.088 0.648 2.16 0.8 ;
        RECT 2.016 0.424 2.088 0.72 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.424 1.872 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.424 1.656 0.72 ;
        RECT 1.512 0.648 1.584 0.8 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.396 1.008 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.72 ;
        RECT 1.08 0.648 1.152 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.424 1.44 0.8 ;
    END
  END B3
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.8 ;
        RECT 0.648 0.728 0.72 0.88 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.9 0.576 0.972 ;
        RECT 0.504 0.28 0.576 0.972 ;
        RECT 0.428 0.28 0.576 0.352 ;
    END
  END C2
  PIN C3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.288 0.576 ;
        RECT 0.072 0.9 0.22 0.972 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END C3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.804 0.9 2.304 0.972 ;
        RECT 2.232 0.252 2.304 0.972 ;
        RECT 1.672 0.252 2.304 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.044 0.252 1.548 0.324 ;
      RECT 1.476 0.108 1.548 0.324 ;
      RECT 1.476 0.108 2.06 0.18 ;
      RECT 0.396 0.108 1.352 0.18 ;
  END
END OAI333_xp33_75t

MACRO OAI33_xp33_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33_xp33_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.8 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.72 ;
        RECT 1.08 0.648 1.152 0.8 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.508 0.728 1.656 0.8 ;
        RECT 1.584 0.28 1.656 0.8 ;
        RECT 1.44 0.504 1.656 0.576 ;
        RECT 1.508 0.28 1.656 0.352 ;
    END
  END A3
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.448 0.792 0.72 ;
        RECT 0.648 0.648 0.72 0.8 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.8 ;
    END
  END B2
  PIN B3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.424 0.36 0.72 ;
        RECT 0.216 0.648 0.288 0.8 ;
    END
  END B3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 1.568 0.972 ;
        RECT 0.072 0.252 0.704 0.324 ;
        RECT 0.072 0.252 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.108 1.444 0.18 ;
  END
END OAI33_xp33_75t

MACRO OR2_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_x1_75t 0 0 ;
  SIZE 1.08 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.944 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.748 ;
        RECT 0.648 0.676 0.72 0.94 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.08 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.08 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.252 0.972 ;
        RECT 0.072 0.108 0.252 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.828 0.872 1.008 0.944 ;
      RECT 0.936 0.108 1.008 0.944 ;
      RECT 0.28 0.504 0.424 0.576 ;
      RECT 0.352 0.108 0.424 0.576 ;
      RECT 0.352 0.108 1.008 0.18 ;
  END
END OR2_x1_75t

MACRO OR2_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_x2_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.728 0.22 0.8 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.9 1.152 0.972 ;
        RECT 1.08 0.108 1.152 0.972 ;
        RECT 0.828 0.108 1.152 0.18 ;
        RECT 0.828 0.736 0.9 0.972 ;
        RECT 0.828 0.108 0.9 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.744 0.972 ;
      RECT 0.672 0.108 0.744 0.972 ;
      RECT 0.672 0.504 0.908 0.576 ;
      RECT 0.376 0.108 0.744 0.18 ;
  END
END OR2_x2_75t

MACRO OR2_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_x4_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.308 0.576 ;
        RECT 0.072 0.728 0.22 0.8 ;
        RECT 0.072 0.108 0.22 0.18 ;
        RECT 0.072 0.108 0.144 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 0.828 0.108 1.656 0.18 ;
        RECT 1.26 0.736 1.332 0.972 ;
        RECT 1.26 0.108 1.332 0.344 ;
        RECT 0.828 0.736 0.9 0.972 ;
        RECT 0.828 0.108 0.9 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.748 0.972 ;
      RECT 0.676 0.108 0.748 0.972 ;
      RECT 0.676 0.504 0.908 0.576 ;
      RECT 0.376 0.108 0.748 0.18 ;
  END
END OR2_x4_75t

MACRO OR2_x6_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_x6_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.252 0.576 0.488 ;
        RECT 0.072 0.252 0.576 0.324 ;
        RECT 0.072 0.252 0.144 0.944 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.612 1.008 0.684 ;
        RECT 0.936 0.424 1.008 0.684 ;
        RECT 0.288 0.424 0.36 0.944 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.9 2.52 0.972 ;
        RECT 2.448 0.108 2.52 0.972 ;
        RECT 1.24 0.108 2.52 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.592 0.756 1.44 0.828 ;
      RECT 1.368 0.28 1.44 0.828 ;
      RECT 1.044 0.28 1.44 0.352 ;
      RECT 1.044 0.108 1.116 0.352 ;
      RECT 0.376 0.108 1.116 0.18 ;
  END
END OR2_x6_75t

MACRO OR3_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_x1_75t 0 0 ;
  SIZE 1.296 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.28 0.364 0.352 ;
        RECT 0.216 0.28 0.288 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.944 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.36 0.792 0.944 ;
        RECT 0.648 0.28 0.72 0.432 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.296 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.296 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.804 1.224 0.876 ;
        RECT 1.152 0.304 1.224 0.876 ;
        RECT 1.044 0.304 1.224 0.376 ;
        RECT 1.044 0.136 1.116 0.376 ;
        RECT 0.936 0.804 1.008 0.944 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 0.292 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.864 0.504 1.008 0.576 ;
      RECT 0.864 0.108 0.936 0.576 ;
      RECT 0.072 0.108 0.936 0.18 ;
  END
END OR3_x1_75t

MACRO OR3_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_x2_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.288 0.576 ;
        RECT 0.072 0.728 0.22 0.8 ;
        RECT 0.072 0.28 0.22 0.352 ;
        RECT 0.072 0.28 0.144 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.72 ;
        RECT 0.648 0.648 0.72 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.732 1.296 0.804 ;
        RECT 1.224 0.304 1.296 0.804 ;
        RECT 1.044 0.304 1.296 0.376 ;
        RECT 1.044 0.732 1.116 0.94 ;
        RECT 1.044 0.136 1.116 0.376 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.936 0.972 ;
      RECT 0.864 0.108 0.936 0.972 ;
      RECT 0.864 0.504 1.048 0.576 ;
      RECT 0.16 0.108 0.936 0.18 ;
  END
END OR3_x2_75t

MACRO OR3_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_x4_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.504 0.288 0.576 ;
        RECT 0.072 0.728 0.22 0.8 ;
        RECT 0.072 0.28 0.22 0.352 ;
        RECT 0.072 0.28 0.144 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.428 0.728 0.576 0.8 ;
        RECT 0.504 0.28 0.576 0.8 ;
        RECT 0.428 0.28 0.576 0.352 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.72 ;
        RECT 0.648 0.648 0.72 0.8 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.044 0.108 1.872 0.18 ;
        RECT 1.476 0.736 1.548 0.972 ;
        RECT 1.476 0.108 1.548 0.344 ;
        RECT 1.044 0.736 1.116 0.972 ;
        RECT 1.044 0.108 1.116 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.16 0.9 0.964 0.972 ;
      RECT 0.892 0.108 0.964 0.972 ;
      RECT 0.892 0.504 1.136 0.576 ;
      RECT 0.16 0.108 0.964 0.18 ;
  END
END OR3_x4_75t

MACRO OR4_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4_x1_75t 0 0 ;
  SIZE 1.512 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.784 ;
        RECT 1.08 0.712 1.152 0.944 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.944 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.864 ;
        RECT 0.648 0.792 0.72 0.944 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.424 0.576 0.944 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.512 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.512 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.272 0.972 ;
        RECT 0.072 0.108 0.272 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.264 0.864 1.44 0.936 ;
      RECT 1.368 0.108 1.44 0.936 ;
      RECT 0.288 0.264 0.36 0.608 ;
      RECT 0.288 0.264 0.468 0.336 ;
      RECT 0.396 0.108 0.468 0.336 ;
      RECT 0.396 0.108 1.44 0.18 ;
  END
END OR4_x1_75t

MACRO OR4_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4_x2_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.364 0.728 1.512 0.8 ;
        RECT 1.44 0.28 1.512 0.8 ;
        RECT 1.364 0.28 1.512 0.352 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.28 1.224 0.864 ;
        RECT 1.08 0.792 1.152 0.944 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.756 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.792 0.792 0.864 0.944 ;
        RECT 0.72 0.424 0.792 0.864 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.9 0.488 0.972 ;
        RECT 0.072 0.108 0.488 0.18 ;
        RECT 0.072 0.108 0.144 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.456 0.9 1.656 0.972 ;
      RECT 1.584 0.108 1.656 0.972 ;
      RECT 0.504 0.264 0.576 0.608 ;
      RECT 0.504 0.264 0.684 0.336 ;
      RECT 0.612 0.108 0.684 0.336 ;
      RECT 0.612 0.108 1.656 0.18 ;
  END
END OR4_x2_75t

MACRO OR4_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4_x4_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.28 1.872 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.28 1.656 0.864 ;
        RECT 1.512 0.792 1.584 0.944 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.28 1.44 0.756 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.224 0.792 1.296 0.944 ;
        RECT 1.152 0.424 1.224 0.864 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.92 0.972 ;
        RECT 0.376 0.108 0.92 0.18 ;
        RECT 0.648 0.108 0.72 0.972 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 1.888 0.9 2.088 0.972 ;
      RECT 2.016 0.108 2.088 0.972 ;
      RECT 0.936 0.264 1.008 0.608 ;
      RECT 0.936 0.264 1.116 0.336 ;
      RECT 1.044 0.108 1.116 0.336 ;
      RECT 1.044 0.108 2.088 0.18 ;
  END
END OR4_x4_75t

MACRO OR5_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5_x1_75t 0 0 ;
  SIZE 1.728 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.716 0.432 0.888 ;
        RECT 0.288 0.28 0.36 0.82 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.9 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.864 ;
        RECT 0.648 0.792 0.72 0.944 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.936 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.86 ;
        RECT 1.08 0.788 1.152 0.94 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.728 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.728 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.4 0.9 1.656 0.972 ;
        RECT 1.584 0.108 1.656 0.972 ;
        RECT 1.396 0.108 1.656 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 0.252 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 1.368 0.252 1.44 0.616 ;
      RECT 1.152 0.252 1.44 0.324 ;
      RECT 1.152 0.108 1.224 0.324 ;
      RECT 0.072 0.108 1.224 0.18 ;
  END
END OR5_x1_75t

MACRO OR5_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5_x2_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.712 0.432 0.888 ;
        RECT 0.288 0.28 0.36 0.82 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.94 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.864 ;
        RECT 0.648 0.792 0.72 0.944 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.936 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.864 ;
        RECT 1.08 0.792 1.152 0.944 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.372 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 0.28 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 1.368 0.252 1.44 0.616 ;
      RECT 1.152 0.252 1.44 0.324 ;
      RECT 1.152 0.108 1.224 0.324 ;
      RECT 0.072 0.108 1.224 0.18 ;
  END
END OR5_x2_75t

MACRO OR5_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR5_x4_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.36 0.668 0.432 0.864 ;
        RECT 0.288 0.28 0.36 0.74 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.94 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.72 0.28 0.792 0.808 ;
        RECT 0.648 0.736 0.72 0.944 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.936 0.28 1.008 0.94 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.152 0.424 1.224 0.796 ;
        RECT 1.08 0.724 1.152 0.944 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.456 0.9 2.304 0.972 ;
        RECT 2.232 0.108 2.304 0.972 ;
        RECT 1.348 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 0.28 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 1.368 0.252 1.44 0.616 ;
      RECT 1.152 0.252 1.44 0.324 ;
      RECT 1.152 0.108 1.224 0.324 ;
      RECT 0.072 0.108 1.224 0.18 ;
  END
END OR5_x4_75t

MACRO SDFH_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFH_x1_75t 0 0 ;
  SIZE 5.4 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.324 0.468 0.396 ;
        RECT 0.396 0.136 0.468 0.396 ;
        RECT 0.216 0.324 0.288 0.8 ;
    END
  END CLK
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.128 0.9 5.328 0.972 ;
        RECT 5.256 0.108 5.328 0.972 ;
        RECT 5.128 0.108 5.328 0.18 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.4 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.4 0.036 ;
    END
  END VSS
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.136 0.432 1.744 0.504 ;
      LAYER M1 ;
        RECT 1.584 0.424 1.656 0.656 ;
      LAYER V1 ;
        RECT 1.584 0.432 1.656 0.504 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.844 0.144 4.916 0.216 ;
      LAYER M1 ;
        RECT 4.824 0.108 5 0.18 ;
        RECT 4.824 0.108 4.896 0.8 ;
        RECT 0.864 0.504 1.244 0.576 ;
        RECT 0.864 0.108 1.032 0.18 ;
        RECT 0.864 0.108 0.936 0.576 ;
      LAYER V1 ;
        RECT 0.864 0.144 0.936 0.216 ;
        RECT 4.824 0.144 4.896 0.216 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.868 0.432 2.36 0.504 ;
      LAYER M1 ;
        RECT 1.94 0.756 2.088 0.828 ;
        RECT 2.016 0.424 2.088 0.828 ;
        RECT 1.844 0.504 2.088 0.576 ;
      LAYER V1 ;
        RECT 2.016 0.432 2.088 0.504 ;
    END
  END SI
  OBS
    LAYER M1 ;
      RECT 4.608 0.9 4.808 0.972 ;
      RECT 4.608 0.136 4.68 0.972 ;
      RECT 4.264 0.9 4.464 0.972 ;
      RECT 4.392 0.108 4.464 0.972 ;
      RECT 3.96 0.108 4.032 0.476 ;
      RECT 3.96 0.108 4.464 0.18 ;
      RECT 3.616 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.744 0.612 4.248 0.684 ;
      RECT 4.176 0.468 4.248 0.684 ;
      RECT 3.4 0.108 3.816 0.18 ;
      RECT 3.168 0.9 3.384 0.972 ;
      RECT 3.312 0.324 3.384 0.972 ;
      RECT 2.88 0.324 3.384 0.396 ;
      RECT 3.204 0.18 3.276 0.396 ;
      RECT 2.88 0.248 2.952 0.396 ;
      RECT 2.32 0.9 2.808 0.972 ;
      RECT 2.736 0.108 2.808 0.972 ;
      RECT 2.736 0.488 3.188 0.56 ;
      RECT 2.536 0.108 2.808 0.18 ;
      RECT 2.448 0.612 2.596 0.684 ;
      RECT 2.448 0.424 2.52 0.684 ;
      RECT 2.232 0.756 2.38 0.828 ;
      RECT 2.232 0.424 2.304 0.828 ;
      RECT 1.044 0.324 1.224 0.396 ;
      RECT 1.152 0.108 1.224 0.396 ;
      RECT 1.152 0.108 2 0.18 ;
      RECT 1.368 0.252 1.44 0.656 ;
      RECT 1.368 0.252 1.516 0.324 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.072 0.9 0.3 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 0.072 0.108 0.272 0.18 ;
      RECT 5.04 0.36 5.112 0.8 ;
      RECT 3.528 0.404 3.6 0.668 ;
      RECT 2.88 0.66 2.952 0.828 ;
      RECT 1.672 0.252 2.436 0.324 ;
      RECT 1.02 0.9 2 0.972 ;
      RECT 1.236 0.756 1.788 0.828 ;
      RECT 0.504 0.484 0.576 0.668 ;
    LAYER M2 ;
      RECT 3.744 0.576 5.132 0.648 ;
      RECT 1.348 0.288 4.7 0.36 ;
      RECT 0.052 0.576 3.6 0.648 ;
      RECT 0.7 0.72 2.972 0.792 ;
    LAYER V1 ;
      RECT 5.04 0.576 5.112 0.648 ;
      RECT 4.608 0.288 4.68 0.36 ;
      RECT 3.744 0.576 3.816 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.88 0.72 2.952 0.792 ;
      RECT 2.448 0.576 2.52 0.648 ;
      RECT 2.232 0.72 2.304 0.792 ;
      RECT 1.368 0.288 1.44 0.36 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.504 0.576 0.576 0.648 ;
      RECT 0.072 0.576 0.144 0.648 ;
  END
END SDFH_x1_75t

MACRO SDFH_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFH_x2_75t 0 0 ;
  SIZE 5.616 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.324 0.468 0.396 ;
        RECT 0.396 0.136 0.468 0.396 ;
        RECT 0.216 0.324 0.288 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.396 1.732 0.468 ;
        RECT 1.584 0.396 1.656 0.656 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.128 0.9 5.472 0.972 ;
        RECT 5.4 0.108 5.472 0.972 ;
        RECT 5.128 0.108 5.472 0.18 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.844 0.144 4.916 0.216 ;
      LAYER M1 ;
        RECT 4.824 0.108 5 0.18 ;
        RECT 4.824 0.108 4.896 0.8 ;
        RECT 1.224 0.504 1.296 0.656 ;
        RECT 0.864 0.504 1.296 0.576 ;
        RECT 0.864 0.108 1.032 0.18 ;
        RECT 0.864 0.108 0.936 0.576 ;
      LAYER V1 ;
        RECT 0.864 0.144 0.936 0.216 ;
        RECT 4.824 0.144 4.896 0.216 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.944 0.424 2.016 0.8 ;
        RECT 1.844 0.504 2.016 0.576 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.616 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.616 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.608 0.9 4.808 0.972 ;
      RECT 4.608 0.136 4.68 0.972 ;
      RECT 4.264 0.9 4.464 0.972 ;
      RECT 4.392 0.108 4.464 0.972 ;
      RECT 3.96 0.108 4.032 0.476 ;
      RECT 3.96 0.108 4.464 0.18 ;
      RECT 3.616 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.744 0.612 4.248 0.684 ;
      RECT 4.176 0.468 4.248 0.684 ;
      RECT 3.4 0.108 3.816 0.18 ;
      RECT 3.168 0.9 3.384 0.972 ;
      RECT 3.312 0.324 3.384 0.972 ;
      RECT 2.88 0.324 3.384 0.396 ;
      RECT 3.204 0.18 3.276 0.396 ;
      RECT 2.88 0.248 2.952 0.396 ;
      RECT 2.32 0.9 2.808 0.972 ;
      RECT 2.736 0.108 2.808 0.972 ;
      RECT 2.736 0.488 3.168 0.56 ;
      RECT 2.536 0.108 2.808 0.18 ;
      RECT 2.448 0.612 2.596 0.684 ;
      RECT 2.448 0.424 2.52 0.684 ;
      RECT 2.232 0.756 2.38 0.828 ;
      RECT 2.232 0.424 2.304 0.828 ;
      RECT 1.044 0.324 1.224 0.396 ;
      RECT 1.152 0.108 1.224 0.396 ;
      RECT 1.152 0.108 2 0.18 ;
      RECT 1.368 0.252 1.44 0.656 ;
      RECT 1.368 0.252 1.516 0.324 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 5.04 0.36 5.112 0.8 ;
      RECT 3.528 0.404 3.6 0.668 ;
      RECT 2.88 0.66 2.952 0.828 ;
      RECT 1.672 0.252 2.436 0.324 ;
      RECT 1.02 0.9 2.024 0.972 ;
      RECT 1.216 0.756 1.788 0.828 ;
      RECT 0.504 0.484 0.576 0.668 ;
    LAYER M2 ;
      RECT 3.744 0.576 5.132 0.648 ;
      RECT 1.348 0.288 4.7 0.36 ;
      RECT 0.036 0.576 3.6 0.648 ;
      RECT 0.7 0.72 2.972 0.792 ;
    LAYER V1 ;
      RECT 5.04 0.576 5.112 0.648 ;
      RECT 4.608 0.288 4.68 0.36 ;
      RECT 3.744 0.576 3.816 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.88 0.72 2.952 0.792 ;
      RECT 2.448 0.576 2.52 0.648 ;
      RECT 2.232 0.72 2.304 0.792 ;
      RECT 1.368 0.288 1.44 0.36 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.504 0.576 0.576 0.648 ;
      RECT 0.036 0.576 0.108 0.648 ;
  END
END SDFH_x2_75t

MACRO SDFH_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFH_x3_75t 0 0 ;
  SIZE 5.832 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.324 0.468 0.396 ;
        RECT 0.396 0.136 0.468 0.396 ;
        RECT 0.288 0.324 0.36 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.396 1.732 0.468 ;
        RECT 1.584 0.396 1.656 0.656 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.128 0.9 5.76 0.972 ;
        RECT 5.688 0.108 5.76 0.972 ;
        RECT 5.128 0.108 5.76 0.18 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.844 0.144 4.916 0.216 ;
      LAYER M1 ;
        RECT 4.824 0.108 5 0.18 ;
        RECT 4.824 0.108 4.896 0.8 ;
        RECT 0.864 0.504 1.244 0.576 ;
        RECT 0.864 0.108 1.032 0.18 ;
        RECT 0.864 0.108 0.936 0.576 ;
      LAYER V1 ;
        RECT 0.864 0.144 0.936 0.216 ;
        RECT 4.824 0.144 4.896 0.216 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.94 0.756 2.088 0.828 ;
        RECT 2.016 0.424 2.088 0.828 ;
        RECT 1.844 0.504 2.088 0.576 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.832 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.832 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.608 0.9 4.808 0.972 ;
      RECT 4.608 0.136 4.68 0.972 ;
      RECT 4.264 0.9 4.464 0.972 ;
      RECT 4.392 0.108 4.464 0.972 ;
      RECT 3.96 0.108 4.032 0.476 ;
      RECT 3.96 0.108 4.464 0.18 ;
      RECT 3.616 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.744 0.612 4.248 0.684 ;
      RECT 4.176 0.468 4.248 0.684 ;
      RECT 3.4 0.108 3.816 0.18 ;
      RECT 3.168 0.9 3.384 0.972 ;
      RECT 3.312 0.324 3.384 0.972 ;
      RECT 2.88 0.324 3.384 0.396 ;
      RECT 3.204 0.18 3.276 0.396 ;
      RECT 2.88 0.248 2.952 0.396 ;
      RECT 2.32 0.9 2.808 0.972 ;
      RECT 2.736 0.108 2.808 0.972 ;
      RECT 2.736 0.488 3.168 0.56 ;
      RECT 2.536 0.108 2.808 0.18 ;
      RECT 2.448 0.612 2.596 0.684 ;
      RECT 2.448 0.424 2.52 0.684 ;
      RECT 2.232 0.756 2.38 0.828 ;
      RECT 2.232 0.424 2.304 0.828 ;
      RECT 1.044 0.324 1.224 0.396 ;
      RECT 1.152 0.108 1.224 0.396 ;
      RECT 1.152 0.108 2 0.18 ;
      RECT 1.368 0.252 1.44 0.656 ;
      RECT 1.368 0.252 1.516 0.324 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.576 0.188 0.648 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 5.04 0.36 5.112 0.8 ;
      RECT 3.528 0.404 3.6 0.668 ;
      RECT 2.88 0.66 2.952 0.828 ;
      RECT 1.672 0.252 2.436 0.324 ;
      RECT 1.02 0.9 2 0.972 ;
      RECT 1.236 0.756 1.788 0.828 ;
      RECT 0.504 0.484 0.576 0.668 ;
    LAYER M2 ;
      RECT 3.744 0.576 5.132 0.648 ;
      RECT 1.348 0.288 4.7 0.36 ;
      RECT 0.076 0.576 3.6 0.648 ;
      RECT 0.7 0.72 2.972 0.792 ;
    LAYER V1 ;
      RECT 5.04 0.576 5.112 0.648 ;
      RECT 4.608 0.288 4.68 0.36 ;
      RECT 3.744 0.576 3.816 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.88 0.72 2.952 0.792 ;
      RECT 2.448 0.576 2.52 0.648 ;
      RECT 2.232 0.72 2.304 0.792 ;
      RECT 1.368 0.288 1.44 0.36 ;
      RECT 0.72 0.72 0.792 0.792 ;
      RECT 0.504 0.576 0.576 0.648 ;
      RECT 0.096 0.576 0.168 0.648 ;
  END
END SDFH_x3_75t

MACRO SDFH_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFH_x4_75t 0 0 ;
  SIZE 6.696 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.252 0.436 0.324 ;
        RECT 0.216 0.252 0.288 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.396 1.872 0.656 ;
        RECT 1.512 0.9 1.836 0.972 ;
        RECT 1.512 0.396 1.872 0.468 ;
        RECT 1.512 0.396 1.584 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.776 0.9 6.624 0.972 ;
        RECT 6.548 0.108 6.624 0.972 ;
        RECT 5.776 0.108 6.624 0.18 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.916 0.288 2.324 0.36 ;
      LAYER M1 ;
        RECT 2.232 0.252 2.396 0.324 ;
        RECT 2.232 0.252 2.304 0.656 ;
        RECT 0.936 0.504 1.156 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
      LAYER V1 ;
        RECT 0.936 0.288 1.008 0.36 ;
        RECT 2.232 0.288 2.304 0.36 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.808 0.108 3.068 0.18 ;
        RECT 2.556 0.3 2.88 0.372 ;
        RECT 2.808 0.108 2.88 0.372 ;
        RECT 2.448 0.424 2.628 0.496 ;
        RECT 2.556 0.3 2.628 0.496 ;
        RECT 2.448 0.424 2.52 0.656 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 6.696 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.696 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.236 0.9 5.544 0.972 ;
      RECT 5.472 0.108 5.544 0.972 ;
      RECT 5.472 0.504 5.788 0.576 ;
      RECT 4.968 0.504 5.132 0.576 ;
      RECT 4.968 0.108 5.04 0.576 ;
      RECT 4.452 0.108 5.544 0.18 ;
      RECT 4.824 0.728 5.328 0.8 ;
      RECT 5.256 0.324 5.328 0.8 ;
      RECT 4.824 0.424 4.896 0.8 ;
      RECT 5.148 0.324 5.328 0.396 ;
      RECT 3.528 0.252 3.6 0.656 ;
      RECT 3.528 0.252 3.924 0.324 ;
      RECT 3.204 0.9 3.816 0.972 ;
      RECT 3.744 0.424 3.816 0.972 ;
      RECT 3.204 0.756 3.276 0.972 ;
      RECT 2.952 0.756 3.276 0.828 ;
      RECT 2.952 0.28 3.024 0.828 ;
      RECT 1.24 0.9 1.44 0.972 ;
      RECT 1.368 0.108 1.44 0.972 ;
      RECT 2.016 0.252 2.088 0.656 ;
      RECT 1.368 0.252 2.088 0.324 ;
      RECT 1.24 0.108 1.44 0.18 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.504 0.108 0.792 0.18 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.108 0.36 0.18 ;
      RECT 4.608 0.424 4.68 0.8 ;
      RECT 4.392 0.28 4.464 0.656 ;
      RECT 4.176 0.424 4.248 0.8 ;
      RECT 3.312 0.28 3.384 0.668 ;
      RECT 3.096 0.28 3.168 0.656 ;
      RECT 2.32 0.9 3.08 0.972 ;
      RECT 2.736 0.484 2.808 0.668 ;
      RECT 1.672 0.108 2.648 0.18 ;
      RECT 1.692 0.756 2.648 0.828 ;
      RECT 0.504 0.424 0.576 0.8 ;
    LAYER M2 ;
      RECT 0.036 0.576 4.7 0.648 ;
      RECT 0.7 0.432 4.484 0.504 ;
    LAYER V1 ;
      RECT 4.608 0.576 4.68 0.648 ;
      RECT 4.392 0.432 4.464 0.504 ;
      RECT 4.176 0.576 4.248 0.648 ;
      RECT 3.312 0.576 3.384 0.648 ;
      RECT 3.096 0.432 3.168 0.504 ;
      RECT 2.736 0.576 2.808 0.648 ;
      RECT 0.72 0.432 0.792 0.504 ;
      RECT 0.504 0.576 0.576 0.648 ;
      RECT 0.036 0.576 0.108 0.648 ;
  END
END SDFH_x4_75t

MACRO SDFL_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFL_x1_75t 0 0 ;
  SIZE 5.4 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.324 0.468 0.396 ;
        RECT 0.396 0.136 0.468 0.396 ;
        RECT 0.288 0.324 0.36 0.656 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.396 1.732 0.468 ;
        RECT 1.584 0.396 1.656 0.656 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.128 0.9 5.328 0.972 ;
        RECT 5.256 0.108 5.328 0.972 ;
        RECT 5.128 0.108 5.328 0.18 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.844 0.144 4.916 0.216 ;
      LAYER M1 ;
        RECT 4.824 0.108 5 0.18 ;
        RECT 4.824 0.108 4.896 0.8 ;
        RECT 0.864 0.504 1.244 0.576 ;
        RECT 0.864 0.108 1.032 0.18 ;
        RECT 0.864 0.108 0.936 0.576 ;
      LAYER V1 ;
        RECT 0.864 0.144 0.936 0.216 ;
        RECT 4.824 0.144 4.896 0.216 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.94 0.756 2.088 0.828 ;
        RECT 2.016 0.424 2.088 0.828 ;
        RECT 1.844 0.504 2.088 0.576 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.4 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.4 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.608 0.9 4.808 0.972 ;
      RECT 4.608 0.136 4.68 0.972 ;
      RECT 4.264 0.9 4.464 0.972 ;
      RECT 4.392 0.108 4.464 0.972 ;
      RECT 3.96 0.108 4.032 0.476 ;
      RECT 3.96 0.108 4.464 0.18 ;
      RECT 3.616 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.744 0.612 4.248 0.684 ;
      RECT 4.176 0.468 4.248 0.684 ;
      RECT 3.4 0.108 3.816 0.18 ;
      RECT 3.168 0.9 3.384 0.972 ;
      RECT 3.312 0.324 3.384 0.972 ;
      RECT 2.88 0.324 3.384 0.396 ;
      RECT 3.204 0.18 3.276 0.396 ;
      RECT 2.88 0.248 2.952 0.396 ;
      RECT 2.32 0.9 2.808 0.972 ;
      RECT 2.736 0.108 2.808 0.972 ;
      RECT 2.736 0.488 3.188 0.56 ;
      RECT 2.536 0.108 2.808 0.18 ;
      RECT 2.448 0.612 2.596 0.684 ;
      RECT 2.448 0.424 2.52 0.684 ;
      RECT 2.232 0.756 2.38 0.828 ;
      RECT 2.232 0.424 2.304 0.828 ;
      RECT 1.044 0.324 1.224 0.396 ;
      RECT 1.152 0.108 1.224 0.396 ;
      RECT 1.152 0.108 2 0.18 ;
      RECT 1.368 0.252 1.44 0.656 ;
      RECT 1.368 0.252 1.516 0.324 ;
      RECT 0.504 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.428 0.756 0.576 0.828 ;
      RECT 0.504 0.484 0.576 0.828 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 5.04 0.36 5.112 0.8 ;
      RECT 3.528 0.404 3.6 0.668 ;
      RECT 2.88 0.66 2.952 0.828 ;
      RECT 1.672 0.252 2.436 0.324 ;
      RECT 1.02 0.9 2 0.972 ;
      RECT 1.236 0.756 1.788 0.828 ;
    LAYER M2 ;
      RECT 3.744 0.576 5.132 0.648 ;
      RECT 1.348 0.288 4.7 0.36 ;
      RECT 0.7 0.576 3.6 0.648 ;
      RECT 0.076 0.72 2.972 0.792 ;
    LAYER V1 ;
      RECT 5.04 0.576 5.112 0.648 ;
      RECT 4.608 0.288 4.68 0.36 ;
      RECT 3.744 0.576 3.816 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.88 0.72 2.952 0.792 ;
      RECT 2.448 0.576 2.52 0.648 ;
      RECT 2.232 0.72 2.304 0.792 ;
      RECT 1.368 0.288 1.44 0.36 ;
      RECT 0.72 0.576 0.792 0.648 ;
      RECT 0.504 0.72 0.576 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END SDFL_x1_75t

MACRO SDFL_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFL_x2_75t 0 0 ;
  SIZE 5.616 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.324 0.468 0.396 ;
        RECT 0.396 0.136 0.468 0.396 ;
        RECT 0.288 0.324 0.36 0.656 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.396 1.732 0.468 ;
        RECT 1.584 0.396 1.656 0.656 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.128 0.9 5.544 0.972 ;
        RECT 5.472 0.108 5.544 0.972 ;
        RECT 5.128 0.108 5.544 0.18 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.844 0.144 4.916 0.216 ;
      LAYER M1 ;
        RECT 4.824 0.108 5 0.18 ;
        RECT 4.824 0.108 4.896 0.8 ;
        RECT 0.864 0.504 1.244 0.576 ;
        RECT 0.864 0.108 1.032 0.18 ;
        RECT 0.864 0.108 0.936 0.576 ;
      LAYER V1 ;
        RECT 0.864 0.144 0.936 0.216 ;
        RECT 4.824 0.144 4.896 0.216 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.94 0.756 2.088 0.828 ;
        RECT 2.016 0.424 2.088 0.828 ;
        RECT 1.844 0.504 2.088 0.576 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.616 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.616 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.608 0.9 4.808 0.972 ;
      RECT 4.608 0.136 4.68 0.972 ;
      RECT 4.264 0.9 4.464 0.972 ;
      RECT 4.392 0.108 4.464 0.972 ;
      RECT 3.96 0.108 4.032 0.476 ;
      RECT 3.96 0.108 4.464 0.18 ;
      RECT 3.616 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.744 0.612 4.248 0.684 ;
      RECT 4.176 0.468 4.248 0.684 ;
      RECT 3.4 0.108 3.816 0.18 ;
      RECT 3.168 0.9 3.384 0.972 ;
      RECT 3.312 0.324 3.384 0.972 ;
      RECT 2.88 0.324 3.384 0.396 ;
      RECT 3.204 0.18 3.276 0.396 ;
      RECT 2.88 0.248 2.952 0.396 ;
      RECT 2.32 0.9 2.808 0.972 ;
      RECT 2.736 0.108 2.808 0.972 ;
      RECT 2.736 0.488 3.168 0.56 ;
      RECT 2.536 0.108 2.808 0.18 ;
      RECT 2.448 0.612 2.596 0.684 ;
      RECT 2.448 0.424 2.52 0.684 ;
      RECT 2.232 0.756 2.38 0.828 ;
      RECT 2.232 0.424 2.304 0.828 ;
      RECT 1.044 0.324 1.224 0.396 ;
      RECT 1.152 0.108 1.224 0.396 ;
      RECT 1.152 0.108 2 0.18 ;
      RECT 1.368 0.252 1.44 0.656 ;
      RECT 1.368 0.252 1.516 0.324 ;
      RECT 0.504 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.428 0.756 0.576 0.828 ;
      RECT 0.504 0.484 0.576 0.828 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 5.04 0.36 5.112 0.8 ;
      RECT 3.528 0.404 3.6 0.668 ;
      RECT 2.88 0.66 2.952 0.828 ;
      RECT 1.672 0.252 2.436 0.324 ;
      RECT 1.02 0.9 2 0.972 ;
      RECT 1.236 0.756 1.788 0.828 ;
    LAYER M2 ;
      RECT 3.744 0.576 5.132 0.648 ;
      RECT 1.348 0.288 4.7 0.36 ;
      RECT 0.7 0.576 3.6 0.648 ;
      RECT 0.076 0.72 2.972 0.792 ;
    LAYER V1 ;
      RECT 5.04 0.576 5.112 0.648 ;
      RECT 4.608 0.288 4.68 0.36 ;
      RECT 3.744 0.576 3.816 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.88 0.72 2.952 0.792 ;
      RECT 2.448 0.576 2.52 0.648 ;
      RECT 2.232 0.72 2.304 0.792 ;
      RECT 1.368 0.288 1.44 0.36 ;
      RECT 0.72 0.576 0.792 0.648 ;
      RECT 0.504 0.72 0.576 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END SDFL_x2_75t

MACRO SDFL_x3_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFL_x3_75t 0 0 ;
  SIZE 5.832 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.324 0.468 0.396 ;
        RECT 0.396 0.136 0.468 0.396 ;
        RECT 0.288 0.324 0.36 0.656 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0.396 1.732 0.468 ;
        RECT 1.584 0.396 1.656 0.656 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.128 0.9 5.76 0.972 ;
        RECT 5.688 0.108 5.76 0.972 ;
        RECT 5.128 0.108 5.76 0.18 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.844 0.144 4.916 0.216 ;
      LAYER M1 ;
        RECT 4.824 0.108 5 0.18 ;
        RECT 4.824 0.108 4.896 0.8 ;
        RECT 0.864 0.504 1.244 0.576 ;
        RECT 0.864 0.108 1.032 0.18 ;
        RECT 0.864 0.108 0.936 0.576 ;
      LAYER V1 ;
        RECT 0.864 0.144 0.936 0.216 ;
        RECT 4.824 0.144 4.896 0.216 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.94 0.756 2.088 0.828 ;
        RECT 2.016 0.424 2.088 0.828 ;
        RECT 1.844 0.504 2.088 0.576 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 5.832 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 5.832 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.608 0.9 4.808 0.972 ;
      RECT 4.608 0.136 4.68 0.972 ;
      RECT 4.264 0.9 4.464 0.972 ;
      RECT 4.392 0.108 4.464 0.972 ;
      RECT 3.96 0.108 4.032 0.476 ;
      RECT 3.96 0.108 4.464 0.18 ;
      RECT 3.616 0.9 3.816 0.972 ;
      RECT 3.744 0.108 3.816 0.972 ;
      RECT 3.744 0.612 4.248 0.684 ;
      RECT 4.176 0.468 4.248 0.684 ;
      RECT 3.4 0.108 3.816 0.18 ;
      RECT 3.168 0.9 3.384 0.972 ;
      RECT 3.312 0.324 3.384 0.972 ;
      RECT 2.88 0.324 3.384 0.396 ;
      RECT 3.204 0.18 3.276 0.396 ;
      RECT 2.88 0.248 2.952 0.396 ;
      RECT 2.32 0.9 2.808 0.972 ;
      RECT 2.736 0.108 2.808 0.972 ;
      RECT 2.736 0.488 3.168 0.56 ;
      RECT 2.536 0.108 2.808 0.18 ;
      RECT 2.448 0.612 2.596 0.684 ;
      RECT 2.448 0.424 2.52 0.684 ;
      RECT 2.232 0.756 2.38 0.828 ;
      RECT 2.232 0.424 2.304 0.828 ;
      RECT 1.044 0.324 1.224 0.396 ;
      RECT 1.152 0.108 1.224 0.396 ;
      RECT 1.152 0.108 2 0.18 ;
      RECT 1.368 0.252 1.44 0.656 ;
      RECT 1.368 0.252 1.516 0.324 ;
      RECT 0.504 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.592 0.108 0.792 0.18 ;
      RECT 0.428 0.756 0.576 0.828 ;
      RECT 0.504 0.484 0.576 0.828 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.72 0.188 0.792 ;
      RECT 0.036 0.108 0.272 0.18 ;
      RECT 5.04 0.36 5.112 0.8 ;
      RECT 3.528 0.404 3.6 0.668 ;
      RECT 2.88 0.66 2.952 0.828 ;
      RECT 1.672 0.252 2.436 0.324 ;
      RECT 1.02 0.9 2 0.972 ;
      RECT 1.236 0.756 1.788 0.828 ;
    LAYER M2 ;
      RECT 3.744 0.576 5.132 0.648 ;
      RECT 1.348 0.288 4.7 0.36 ;
      RECT 0.7 0.576 3.6 0.648 ;
      RECT 0.076 0.72 2.972 0.792 ;
    LAYER V1 ;
      RECT 5.04 0.576 5.112 0.648 ;
      RECT 4.608 0.288 4.68 0.36 ;
      RECT 3.744 0.576 3.816 0.648 ;
      RECT 3.528 0.576 3.6 0.648 ;
      RECT 2.88 0.72 2.952 0.792 ;
      RECT 2.448 0.576 2.52 0.648 ;
      RECT 2.232 0.72 2.304 0.792 ;
      RECT 1.368 0.288 1.44 0.36 ;
      RECT 0.72 0.576 0.792 0.648 ;
      RECT 0.504 0.72 0.576 0.792 ;
      RECT 0.096 0.72 0.168 0.792 ;
  END
END SDFL_x3_75t

MACRO SDFL_x4_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFL_x4_75t 0 0 ;
  SIZE 6.696 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.216 0.252 0.436 0.324 ;
        RECT 0.216 0.252 0.288 0.8 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.8 0.396 1.872 0.656 ;
        RECT 1.512 0.9 1.836 0.972 ;
        RECT 1.512 0.396 1.872 0.468 ;
        RECT 1.512 0.396 1.584 0.972 ;
    END
  END D
  PIN QN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 5.776 0.9 6.624 0.972 ;
        RECT 6.548 0.108 6.624 0.972 ;
        RECT 5.776 0.108 6.624 0.18 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.916 0.288 2.324 0.36 ;
      LAYER M1 ;
        RECT 2.232 0.252 2.396 0.324 ;
        RECT 2.232 0.252 2.304 0.656 ;
        RECT 0.936 0.504 1.156 0.576 ;
        RECT 0.936 0.9 1.084 0.972 ;
        RECT 0.936 0.108 1.084 0.18 ;
        RECT 0.936 0.108 1.008 0.972 ;
      LAYER V1 ;
        RECT 0.936 0.288 1.008 0.36 ;
        RECT 2.232 0.288 2.304 0.36 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.808 0.108 3.068 0.18 ;
        RECT 2.556 0.3 2.88 0.372 ;
        RECT 2.808 0.108 2.88 0.372 ;
        RECT 2.448 0.424 2.628 0.496 ;
        RECT 2.556 0.3 2.628 0.496 ;
        RECT 2.448 0.424 2.52 0.656 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 6.696 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 6.696 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 4.236 0.9 5.544 0.972 ;
      RECT 5.472 0.108 5.544 0.972 ;
      RECT 5.472 0.504 5.788 0.576 ;
      RECT 4.968 0.504 5.132 0.576 ;
      RECT 4.968 0.108 5.04 0.576 ;
      RECT 4.452 0.108 5.544 0.18 ;
      RECT 4.824 0.728 5.328 0.8 ;
      RECT 5.256 0.324 5.328 0.8 ;
      RECT 4.824 0.424 4.896 0.8 ;
      RECT 5.148 0.324 5.328 0.396 ;
      RECT 3.528 0.252 3.6 0.656 ;
      RECT 3.528 0.252 3.924 0.324 ;
      RECT 3.204 0.9 3.816 0.972 ;
      RECT 3.744 0.424 3.816 0.972 ;
      RECT 3.204 0.756 3.276 0.972 ;
      RECT 2.952 0.756 3.276 0.828 ;
      RECT 2.952 0.28 3.024 0.828 ;
      RECT 1.24 0.9 1.44 0.972 ;
      RECT 1.368 0.108 1.44 0.972 ;
      RECT 2.016 0.252 2.088 0.656 ;
      RECT 1.368 0.252 2.088 0.324 ;
      RECT 1.24 0.108 1.44 0.18 ;
      RECT 0.592 0.9 0.792 0.972 ;
      RECT 0.72 0.108 0.792 0.972 ;
      RECT 0.504 0.108 0.792 0.18 ;
      RECT 0.036 0.9 0.272 0.972 ;
      RECT 0.036 0.108 0.108 0.972 ;
      RECT 0.036 0.108 0.36 0.18 ;
      RECT 4.608 0.424 4.68 0.8 ;
      RECT 4.392 0.28 4.464 0.656 ;
      RECT 4.176 0.424 4.248 0.8 ;
      RECT 3.312 0.28 3.384 0.668 ;
      RECT 3.096 0.28 3.168 0.656 ;
      RECT 2.32 0.9 3.08 0.972 ;
      RECT 2.736 0.484 2.808 0.668 ;
      RECT 1.672 0.108 2.648 0.18 ;
      RECT 1.692 0.756 2.648 0.828 ;
      RECT 0.504 0.412 0.576 0.8 ;
    LAYER M2 ;
      RECT 0.7 0.576 4.7 0.648 ;
      RECT 0.036 0.432 4.484 0.504 ;
    LAYER V1 ;
      RECT 4.608 0.576 4.68 0.648 ;
      RECT 4.392 0.432 4.464 0.504 ;
      RECT 4.176 0.576 4.248 0.648 ;
      RECT 3.312 0.576 3.384 0.648 ;
      RECT 3.096 0.432 3.168 0.504 ;
      RECT 2.736 0.576 2.808 0.648 ;
      RECT 0.72 0.576 0.792 0.648 ;
      RECT 0.504 0.432 0.576 0.504 ;
      RECT 0.036 0.432 0.108 0.504 ;
  END
END SDFL_x4_75t

MACRO TAPCELL_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TAPCELL_75t 0 0 ;
  SIZE 0.432 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.432 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.432 0.036 ;
    END
  END VSS
END TAPCELL_75t

MACRO TAPCELL_WITH_FILLER_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TAPCELL_WITH_FILLER_75t 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
END TAPCELL_WITH_FILLER_75t

MACRO TIEHI_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHI_x1_75t 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN H
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.376 0.9 0.576 0.972 ;
        RECT 0.504 0.28 0.576 0.972 ;
        RECT 0.268 0.28 0.576 0.352 ;
    END
  END H
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.072 0.512 0.38 0.584 ;
      RECT 0.072 0.108 0.144 0.584 ;
      RECT 0.072 0.108 0.272 0.18 ;
  END
END TIEHI_x1_75t

MACRO TIELO_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELO_x1_75t 0 0 ;
  SIZE 0.648 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN L
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.268 0.728 0.576 0.8 ;
        RECT 0.504 0.108 0.576 0.8 ;
        RECT 0.376 0.108 0.576 0.18 ;
    END
  END L
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 0.648 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 0.648 0.036 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 0.272 0.972 ;
      RECT 0.072 0.496 0.144 0.972 ;
      RECT 0.072 0.496 0.38 0.568 ;
  END
END TIELO_x1_75t

MACRO XNOR2_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_x1_75t 0 0 ;
  SIZE 2.16 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.16 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.16 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.9 1.568 0.972 ;
        RECT 1.368 0.268 1.568 0.34 ;
        RECT 1.368 0.268 1.44 0.972 ;
        RECT 0.808 0.748 1.44 0.82 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.484 0.288 1.976 0.36 ;
      LAYER M1 ;
        RECT 1.8 0.288 1.976 0.36 ;
        RECT 1.8 0.288 1.872 0.596 ;
        RECT 1.152 0.288 1.224 0.648 ;
        RECT 1.048 0.288 1.224 0.36 ;
        RECT 0.504 0.268 0.576 0.688 ;
      LAYER V1 ;
        RECT 0.504 0.288 0.576 0.36 ;
        RECT 1.068 0.288 1.14 0.36 ;
        RECT 1.884 0.288 1.956 0.36 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.268 0.432 0.812 0.504 ;
      LAYER M1 ;
        RECT 0.72 0.336 0.792 0.66 ;
        RECT 0.288 0.268 0.36 0.596 ;
      LAYER V1 ;
        RECT 0.288 0.432 0.36 0.504 ;
        RECT 0.72 0.432 0.792 0.504 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 1.584 0.72 2 0.792 ;
      RECT 1.584 0.428 1.656 0.792 ;
      RECT 0.072 0.72 0.272 0.792 ;
      RECT 0.072 0.108 0.144 0.792 ;
      RECT 0.072 0.108 0.272 0.18 ;
      RECT 0.808 0.108 1.784 0.18 ;
      RECT 0.592 0.9 1.136 0.972 ;
    LAYER M2 ;
      RECT 0.16 0.72 2 0.792 ;
    LAYER V1 ;
      RECT 1.908 0.72 1.98 0.792 ;
      RECT 0.18 0.72 0.252 0.792 ;
  END
END XNOR2_x1_75t

MACRO XNOR2_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_x2_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.044 0.9 1.76 0.972 ;
        RECT 1.688 0.504 1.76 0.972 ;
        RECT 1.564 0.504 1.76 0.576 ;
        RECT 1.044 0.732 1.116 0.972 ;
        RECT 0.504 0.732 1.116 0.804 ;
        RECT 0.504 0.424 0.576 0.804 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.756 1.588 0.828 ;
        RECT 1.368 0.424 1.44 0.828 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.888 0.9 2.304 0.972 ;
        RECT 2.232 0.108 2.304 0.972 ;
        RECT 1.888 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 0.252 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 1.908 0.252 1.98 0.604 ;
      RECT 1.692 0.252 1.98 0.324 ;
      RECT 1.692 0.108 1.764 0.324 ;
      RECT 0.072 0.108 1.764 0.18 ;
      RECT 1.208 0.252 1.28 0.78 ;
      RECT 0.288 0.252 0.36 0.596 ;
      RECT 0.288 0.252 1.568 0.324 ;
      RECT 0.396 0.9 0.92 0.972 ;
  END
END XNOR2_x2_75t

MACRO XNOR2_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_xp5_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.252 1.44 0.656 ;
        RECT 0.828 0.252 1.44 0.324 ;
        RECT 0.828 0.108 0.9 0.324 ;
        RECT 0.216 0.108 0.9 0.18 ;
        RECT 0.216 0.108 0.288 0.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.28 0.576 0.8 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.692 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.376 0.9 0.72 0.972 ;
      RECT 0.648 0.3 0.72 0.972 ;
      RECT 0.648 0.756 1.656 0.828 ;
      RECT 1.584 0.484 1.656 0.828 ;
      RECT 1.044 0.108 1.548 0.18 ;
  END
END XNOR2_xp5_75t

MACRO XOR2_x1_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_x1_75t 0 0 ;
  SIZE 2.592 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 1.192 0.72 2.108 0.792 ;
      LAYER M1 ;
        RECT 2.016 0.472 2.088 0.8 ;
        RECT 1.22 0.504 1.46 0.576 ;
        RECT 0.852 0.74 1.292 0.812 ;
        RECT 1.22 0.504 1.292 0.812 ;
        RECT 0.072 0.9 0.924 0.972 ;
        RECT 0.852 0.74 0.924 0.972 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.136 0.144 0.972 ;
      LAYER V1 ;
        RECT 1.22 0.72 1.292 0.792 ;
        RECT 2.016 0.72 2.088 0.792 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.592 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.592 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.024 0.108 2.448 0.18 ;
        RECT 1.672 0.7 1.872 0.772 ;
        RECT 1.8 0.108 1.872 0.772 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.484 0.288 2.324 0.36 ;
      LAYER M1 ;
        RECT 2.232 0.252 2.304 0.596 ;
        RECT 2.104 0.252 2.304 0.324 ;
        RECT 0.504 0.252 0.576 0.596 ;
        RECT 0.428 0.252 0.576 0.324 ;
      LAYER V1 ;
        RECT 0.504 0.288 0.576 0.36 ;
        RECT 2.232 0.288 2.304 0.36 ;
    END
  END B
  OBS
    LAYER M1 ;
      RECT 0.696 0.108 0.768 0.752 ;
      RECT 1.584 0.252 1.656 0.596 ;
      RECT 0.696 0.252 1.656 0.324 ;
      RECT 0.696 0.108 0.772 0.324 ;
      RECT 0.368 0.108 0.772 0.18 ;
      RECT 1.024 0.9 2.432 0.972 ;
  END
END XOR2_x1_75t

MACRO XOR2_x2_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_x2_75t 0 0 ;
  SIZE 2.376 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.368 0.252 1.516 0.324 ;
        RECT 1.368 0.252 1.44 0.652 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.688 0.108 1.76 0.652 ;
        RECT 1.564 0.504 1.76 0.576 ;
        RECT 1.044 0.108 1.76 0.18 ;
        RECT 0.504 0.276 1.116 0.348 ;
        RECT 1.044 0.108 1.116 0.348 ;
        RECT 0.504 0.276 0.576 0.6 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 2.376 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 2.376 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.888 0.9 2.304 0.972 ;
        RECT 2.232 0.108 2.304 0.972 ;
        RECT 1.888 0.108 2.304 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.9 1.764 0.972 ;
      RECT 1.692 0.756 1.764 0.972 ;
      RECT 0.072 0.108 0.144 0.972 ;
      RECT 1.692 0.756 1.98 0.828 ;
      RECT 1.908 0.476 1.98 0.828 ;
      RECT 0.072 0.108 0.252 0.18 ;
      RECT 0.288 0.756 1.568 0.828 ;
      RECT 1.208 0.3 1.28 0.828 ;
      RECT 0.288 0.484 0.36 0.828 ;
      RECT 0.396 0.108 0.92 0.18 ;
  END
END XOR2_x2_75t

MACRO XOR2_xp5_75t
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_xp5_75t 0 0 ;
  SIZE 1.944 BY 1.08 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.828 0.756 1.44 0.828 ;
        RECT 1.368 0.48 1.44 0.828 ;
        RECT 0.072 0.9 0.9 0.972 ;
        RECT 0.828 0.756 0.9 0.972 ;
        RECT 0.072 0.504 0.312 0.576 ;
        RECT 0.072 0.136 0.144 0.972 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.424 0.756 0.576 0.828 ;
        RECT 0.504 0.252 0.576 0.828 ;
        RECT 0.428 0.252 0.576 0.324 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 1.044 1.944 1.116 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M1 ;
        RECT 0 -0.036 1.944 0.036 ;
    END
  END VSS
  PIN Y
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.692 0.9 1.872 0.972 ;
        RECT 1.8 0.108 1.872 0.972 ;
        RECT 1.024 0.108 1.872 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.648 0.108 0.72 0.78 ;
      RECT 1.584 0.252 1.656 0.596 ;
      RECT 0.648 0.252 1.656 0.324 ;
      RECT 0.376 0.108 0.72 0.18 ;
      RECT 1.024 0.9 1.548 0.972 ;
  END
END XOR2_xp5_75t

END LIBRARY
